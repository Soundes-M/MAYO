--------------------------------------------------------------------------------
-- Title       : <Title Block>
-- Project     : Default Project Name
--------------------------------------------------------------------------------
-- File        : MAYO_BRAM_Arbiter.vhd
-- Author      : User Name <user.email@user.company.com>
-- Company     : User Company Name
-- Created     : Mon Oct  3 12:33:18 2022
-- Last update : Sat Apr 29 18:37:06 2023
-- Platform    : Default Part Number
-- Standard    : <VHDL-2008 | VHDL-2002 | VHDL-1993 | VHDL-1987>
--------------------------------------------------------------------------------
-- Copyright (c) 2022 User Company Name
-------------------------------------------------------------------------------
-- Description: Pass through for BRAM signals. 
-- Works only in Sign
-- Leave ports open if not needed.
--------------------------------------------------------------------------------
-- Revisions:  Revisions and documentation are controlled by
-- the revision control system (RCS).  The RCS should be consulted
-- on revision history.
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

use work.MAYO_COMMON.all;
use work.UTILS_COMMON.all;

entity mayo_bram_arbiter is
	port (

		-- Sign Main FSM
		BRAM_sign_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_sign_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_sign_en   : in  std_logic;
		BRAM_sign_rst  : in  std_logic;
		BRAM_sign_we   : in  std_logic_vector (3 downto 0);
		BRAM_sign_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		BRAM_add_vec_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_add_vec_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_add_vec_en   : in  std_logic;
		BRAM_add_vec_rst  : in  std_logic;
		BRAM_add_vec_we   : in  std_logic_vector (3 downto 0);
		BRAM_add_vec_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		BRAM_lin_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_lin_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_lin_en   : in  std_logic;
		BRAM_lin_rst  : in  std_logic;
		BRAM_lin_we   : in  std_logic_vector (3 downto 0);
		BRAM_lin_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		BRAM_neg_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_neg_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_neg_en   : in  std_logic;
		BRAM_neg_rst  : in  std_logic;
		BRAM_neg_we   : in  std_logic_vector (3 downto 0);
		BRAM_neg_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		BRAM_red_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_red_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_red_en   : in  std_logic;
		BRAM_red_rst  : in  std_logic;
		BRAM_red_we   : in  std_logic_vector (3 downto 0);
		BRAM_red_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		BRAM_sam_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_sam_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_sam_en   : in  std_logic;
		BRAM_sam_rst  : in  std_logic;
		BRAM_sam_we   : in  std_logic_vector (3 downto 0);
		BRAM_sam_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		BRAM_memcpy0_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_memcpy0_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_memcpy0_en   : in  std_logic;
		BRAM_memcpy0_rst  : in  std_logic;
		BRAM_memcpy0_we   : in  std_logic_vector (3 downto 0);
		BRAM_memcpy0_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		BRAM_memcpy1_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_memcpy1_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_memcpy1_en   : in  std_logic;
		BRAM_memcpy1_rst  : in  std_logic;
		BRAM_memcpy1_we   : in  std_logic_vector (3 downto 0);
		BRAM_memcpy1_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		BRAM_p1p1t_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_p1p1t_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_p1p1t_en   : in  std_logic;
		BRAM_p1p1t_rst  : in  std_logic;
		BRAM_p1p1t_we   : in  std_logic_vector (3 downto 0);
		BRAM_p1p1t_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		BRAM_red_ext_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_red_ext_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_red_ext_en   : in  std_logic;
		BRAM_red_ext_rst  : in  std_logic;
		BRAM_red_ext_we   : in  std_logic_vector (3 downto 0);
		BRAM_red_ext_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		BRAM_sam_vin_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_sam_vin_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_sam_vin_en   : in  std_logic;
		BRAM_sam_vin_rst  : in  std_logic;
		BRAM_sam_vin_we   : in  std_logic_vector (3 downto 0);
		BRAM_sam_vin_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		BRAM_sam_oil_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_sam_oil_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_sam_oil_en   : in  std_logic;
		BRAM_sam_oil_rst  : in  std_logic;
		BRAM_sam_oil_we   : in  std_logic_vector (3 downto 0);
		BRAM_sam_oil_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		BRAM_add_oil_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_add_oil_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_add_oil_en   : in  std_logic;
		BRAM_add_oil_rst  : in  std_logic;
		BRAM_add_oil_we   : in  std_logic_vector (3 downto 0);
		BRAM_add_oil_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		-- Hash 
		BRAM_hash_din  : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_hash_addr : in  std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_hash_en   : in  std_logic;
		BRAM_hash_rst  : in  std_logic;
		BRAM_hash_we   : in  std_logic_vector (3 downto 0);
		BRAM_hash_dout : out std_logic_vector(PORT_WIDTH-1 downto 0);

		-- OUTPUT
		BRAM_din  : out std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_addr : out std_logic_vector(PORT_WIDTH-1 downto 0);
		BRAM_en   : out std_logic;
		BRAM_rst  : out std_logic;
		BRAM_we   : out std_logic_vector (3 downto 0);
		BRAM_dout : in  std_logic_vector(PORT_WIDTH-1 downto 0);

		-- FSM From MAYO Control
		add_vec_control : in std_logic;
		lin_control     : in std_logic;
		neg_control     : in std_logic;
		red_control     : in std_logic;
		sam_control     : in std_logic;
		hash_control    : in std_logic;
		memcpy0_control : in std_logic;
		memcpy1_control : in std_logic;
		p1p1t_control   : in std_logic;
		red_ext_control : in std_logic;
		sam_vin_control : in std_logic;
		sam_oil_control : in std_logic;
		add_oil_control : in std_logic;
		-- Sign control
		bram_control : in std_logic

	);
end entity mayo_bram_arbiter;

architecture Behavioral of mayo_bram_arbiter is

begin
	BRAM_din <= BRAM_sign_din when (bram_control = '1')
	else BRAM_add_vec_din     when (add_vec_control = '1')
	else BRAM_lin_din         when (lin_control = '1')
	else BRAM_neg_din         when (neg_control = '1')
	else BRAM_red_din         when (red_control ='1')
	else BRAM_sam_din         when (sam_control = '1')
	else BRAM_hash_din        when (hash_control = '1')
	else BRAM_memcpy0_din     when (memcpy0_control = '1')
	else BRAM_memcpy1_din     when (memcpy1_control = '1')
	else BRAM_p1p1t_din       when (p1p1t_control = '1')
	else BRAM_red_ext_din     when (red_ext_control = '1')
	else BRAM_sam_vin_din     when (sam_vin_control = '1')
	else BRAM_sam_oil_din     when (sam_oil_control = '1')
	else BRAM_add_oil_din     when (add_oil_control = '1')
	else (others => '0');

	BRAM_addr <= BRAM_sign_addr when (bram_control = '1')
	else BRAM_add_vec_addr      when (add_vec_control = '1')
	else BRAM_lin_addr          when (lin_control = '1')
	else BRAM_neg_addr          when (neg_control = '1')
	else BRAM_red_addr          when (red_control ='1')
	else BRAM_sam_addr          when (sam_control = '1')
	else BRAM_hash_addr         when (hash_control = '1')
	else BRAM_memcpy0_addr      when (memcpy0_control = '1')
	else BRAM_memcpy1_addr      when (memcpy1_control = '1')
	else BRAM_p1p1t_addr        when (p1p1t_control = '1')
	else BRAM_red_ext_addr      when (red_ext_control = '1')
	else BRAM_sam_vin_addr      when (sam_vin_control = '1')
	else BRAM_sam_oil_addr      when (sam_oil_control = '1')
	else BRAM_add_oil_addr      when (add_oil_control = '1')
	else (others => '0');

	BRAM_we <= BRAM_sign_we when (bram_control = '1')
	else BRAM_add_vec_we    when (add_vec_control = '1')
	else BRAM_lin_we        when (lin_control = '1')
	else BRAM_neg_we        when (neg_control = '1')
	else BRAM_red_we        when (red_control ='1')
	else BRAM_sam_we        when (sam_control = '1')
	else BRAM_hash_we       when (hash_control = '1')
	else BRAM_memcpy0_we    when (memcpy0_control = '1')
	else BRAM_memcpy1_we    when (memcpy1_control = '1')
	else BRAM_p1p1t_we      when (p1p1t_control = '1')
	else BRAM_red_ext_we    when (red_ext_control = '1')
	else BRAM_sam_vin_we    when (sam_vin_control = '1')
	else BRAM_sam_oil_we    when (sam_oil_control = '1')
	else BRAM_add_oil_we    when (add_oil_control = '1')
	else (others => '0');

	BRAM_en <= '1' when ( (BRAM_add_vec_en = '1')
			or (BRAM_lin_en = '1')
			or (BRAM_neg_en = '1')
			or (BRAM_red_en = '1')
			or (BRAM_sign_en = '1')
			or (BRAM_sam_en = '1')
			or (BRAM_hash_en = '1')
			or (BRAM_memcpy0_en = '1')
			or (BRAM_memcpy1_en = '1')
			or (BRAM_p1p1t_en = '1')
			or (BRAM_red_ext_en = '1')
			or (BRAM_sam_vin_en = '1')
			or (BRAM_sam_oil_en = '1')
			or (BRAM_add_oil_en = '1'))
	else '0;

	BRAM_rst <= '1' when ( (BRAM_add_vec_rst = '1')
			or (BRAM_lin_rst = '1')
			or (BRAM_neg_rst = '1')
			or (BRAM_red_rst = '1')
			or (BRAM_sign_rst = '1')
			or (BRAM_sam_rst = '1')
			or (BRAM_hash_rst = '1')
			or (BRAM_memcpy0_rst = '1')
			or (BRAM_memcpy1_rst = '1')
			or (BRAM_p1p1t_rst = '1')
			or (BRAM_red_ext_rst = '1')
			or (BRAM_sam_vin_rst = '1')
			or (BRAM_sam_oil_rst = '1')
			or (BRAM_add_oil_rst = '1'))
	else '0';

	BRAM_sign_dout    <= BRAM_dout when (bram_control = '1') else (others    => '0');
	BRAM_add_vec_dout <= BRAM_dout when (add_vec_control = '1') else (others => '0');
	BRAM_lin_dout     <= BRAM_dout when (lin_control = '1') else (others     => '0');
	BRAM_neg_dout     <= BRAM_dout when (neg_control = '1') else (others     => '0');
	BRAM_red_dout     <= BRAM_dout when (red_control = '1') else (others     => '0');
	BRAM_sam_dout     <= BRAM_dout when (sam_control = '1') else (others     => '0');
	BRAM_hash_dout    <= BRAM_dout when (hash_control = '1') else (others    => '0');
	BRAM_memcpy0_dout <= BRAM_dout when (memcpy0_control = '1') else (others => '0');
	BRAM_memcpy1_dout <= BRAM_dout when (memcpy1_control = '1') else (others => '0');
	BRAM_p1p1t_dout   <= BRAM_dout when (p1p1t_control = '1') else (others   => '0');
	BRAM_red_ext_dout <= BRAM_dout when (red_ext_control = '1') else (others => '0');
	BRAM_sam_vin_dout <= BRAM_dout when (sam_vin_control = '1') else (others => '0');
	BRAM_sam_oil_dout <= BRAM_dout when (sam_oil_control = '1') else (others => '0');
	BRAM_add_oil_dout <= BRAM_dout when (add_oil_control = '1') else (others => '0');

end architecture Behavioral;