library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity gsmith_generated is
	port (
		clk      : in  std_logic;
		rst      : in  std_logic;
		enable   : in  std_logic;
		lo       : in  std_logic;
		fet      : in  std_logic;
		data_in  : in  std_logic_vector(7 downto 0);
		data_out : out std_logic_vector(7 downto 0);
		i        : in  std_logic_vector(31 downto 0);
		j        : in  std_logic_vector(31 downto 0);
		done     : out std_logic
	);

end entity gsmith_generated;

architecture behav of gsmith_generated is
	component basic_cell is
		port (
			clk                : in  std_logic;
			rst                : in  std_logic;
			en                 : in  std_logic;
			load               : in  std_logic;
			fetch              : in  std_logic;
			data_in            : in  std_logic_vector(7 downto 0);
			data_out           : out std_logic_vector(7 downto 0);
			out1               : out std_logic_vector(7 downto 0); -- Upper neighbor
			out2               : out std_logic_vector(7 downto 0); -- Upper left
			lock_lower_row_out : out std_logic;                    -- Upper neighbor
			lock_lower_row_in  : in  std_logic;                    -- Lower neighbor
			in1                : in  std_logic_vector(7 downto 0); -- Lower neighbor
			in2                : in  std_logic_vector(7 downto 0); -- Lower right
			lock_row           : in  std_logic;
			piv_found          : in  std_logic;
			row_data           : in  std_logic_vector(7 downto 0);
			col_data           : in  std_logic_vector(7 downto 0)
		);
	end component basic_cell;

	component pivot_cell is
		port (
			clk       : in  std_logic;
			rst       : in  std_logic;
			en        : in  std_logic;
			load      : in  std_logic;
			fetch     : in  std_logic;
			data_in   : in  std_logic_vector(7 downto 0);
			data_out  : out std_logic_vector(7 downto 0);
			in1       : in  std_logic_vector(7 downto 0);
			in2       : in  std_logic_vector(7 downto 0);
			row_data  : out std_logic_vector(7 downto 0);
			piv_found : out std_logic
		);
	end component pivot_cell;

	component pivotRow_cell is
		port (
			clk       : in  std_logic;
			rst       : in  std_logic;
			en        : in  std_logic;
			load      : in  std_logic;
			fetch     : in  std_logic;
			data_in   : in  std_logic_vector(7 downto 0);
			data_out  : out std_logic_vector(7 downto 0);
			out1      : out std_logic_vector(7 downto 0);
			out2      : out std_logic_vector(7 downto 0);
			in1       : in  std_logic_vector(7 downto 0);
			in2       : in  std_logic_vector(7 downto 0);
			piv_found : in  std_logic;
			row_data  : in  std_logic_vector(7 downto 0);
			col_data  : out std_logic_vector(7 downto 0)
		);
	end component pivotRow_cell;

	component pivotCol_cell is
		port (
			clk                : in  std_logic;
			rst                : in  std_logic;
			en                 : in  std_logic;
			load               : in  std_logic;
			fetch              : in  std_logic;
			data_in            : in  std_logic_vector(7 downto 0);
			data_out           : out std_logic_vector(7 downto 0);
			out1               : out std_logic_vector(7 downto 0); -- Upper neighbor
			lock_lower_row_out : out std_logic;                    -- Upper neighbor
			lock_lower_row_in  : in  std_logic;                    -- Lower neighbor
			in1                : in  std_logic_vector(7 downto 0); -- Lower neighbor
			in2                : in  std_logic_vector(7 downto 0); -- Lower right
			lock_row           : in  std_logic;
			piv_found          : in  std_logic;
			row_data           : out std_logic_vector(7 downto 0)
		);
	end component pivotCol_cell;

	-- Matrix Size (ROWS*COLS)
	CONSTANT ROWS : integer := 60;
	CONSTANT COLS : integer := 61;

	signal s_piv_found : std_logic;
	type vector8 is array (natural range <>) of std_logic_vector(7 downto 0);
	type vector8_2d is array (0 to ROWS-1, 0 to COLS-1) of std_logic_vector(7 downto 0);
	type vector1_2d is array (0 to ROWS-1, 0 to COLS-1) of std_logic;
	signal s_row_data : vector8(0 to ROWS-1);
	signal s_col_data : vector8(0 to COLS-1);
	signal s_in1      : vector8_2d;
	signal s_in2      : vector8_2d;
	signal s_out1     : vector8_2d;
	signal s_out2     : vector8_2d;
	signal s_data_in  : vector8_2d;
	signal s_data_out : vector8_2d;
	signal s_fetch    : vector1_2d;
	signal s_load     : vector1_2d;
	signal tmp        : std_logic;
	type vector1 is array (natural range <>) of std_logic;
	signal s_locks_lower_in  : vector1_2d;
	signal s_locks_lower_out : vector1_2d;
	signal s_locks           : vector1(0 to ROWS-1); -- also called 'used' flag
	signal en                : std_logic := '0';
	signal s_i, s_j          : unsigned(31 downto 0);
	function check_locks(locks : vector1) return std_logic is
		variable result            : std_logic := '1';
	begin
		for i in locks'range loop
			if locks(i) = '0' then
				result := '0';
				exit;
			end if;
		end loop;
		return result;
	end function;

begin
		pivot_gen : pivot_cell port map (
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,0),
			fetch     => s_fetch(0,0),
			data_in   => s_data_in(0,0),
			data_out  => s_data_out(0,0),
			in1       => s_in1(0,0),
			in2       => s_in2(0,0),
			row_data  => s_row_data(0),
			piv_found => s_piv_found
		);
	s_in1(0,0) <= s_out1(1,0);
	s_in2(0,0) <= s_out2(1,1);


		--Pivot Rows-----------
		piv_row_1 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,1),
			fetch     => s_fetch(0,1),
			data_in   => s_data_in(0,1),
			data_out  => s_data_out(0,1),
			out1      => s_out1(0,1),
			out2      => s_out2(0,1),
			in1       => s_in1(0,1),
			in2       => s_in2(0,1),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(1)
		);
	s_in1(0,1) <= s_out1(1,1);
	s_in2(0,1) <= s_out2(1,2);

		piv_row_2 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,2),
			fetch     => s_fetch(0,2),
			data_in   => s_data_in(0,2),
			data_out  => s_data_out(0,2),
			out1      => s_out1(0,2),
			out2      => s_out2(0,2),
			in1       => s_in1(0,2),
			in2       => s_in2(0,2),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(2)
		);
	s_in1(0,2) <= s_out1(1,2);
	s_in2(0,2) <= s_out2(1,3);

		piv_row_3 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,3),
			fetch     => s_fetch(0,3),
			data_in   => s_data_in(0,3),
			data_out  => s_data_out(0,3),
			out1      => s_out1(0,3),
			out2      => s_out2(0,3),
			in1       => s_in1(0,3),
			in2       => s_in2(0,3),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(3)
		);
	s_in1(0,3) <= s_out1(1,3);
	s_in2(0,3) <= s_out2(1,4);

		piv_row_4 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,4),
			fetch     => s_fetch(0,4),
			data_in   => s_data_in(0,4),
			data_out  => s_data_out(0,4),
			out1      => s_out1(0,4),
			out2      => s_out2(0,4),
			in1       => s_in1(0,4),
			in2       => s_in2(0,4),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(4)
		);
	s_in1(0,4) <= s_out1(1,4);
	s_in2(0,4) <= s_out2(1,5);

		piv_row_5 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,5),
			fetch     => s_fetch(0,5),
			data_in   => s_data_in(0,5),
			data_out  => s_data_out(0,5),
			out1      => s_out1(0,5),
			out2      => s_out2(0,5),
			in1       => s_in1(0,5),
			in2       => s_in2(0,5),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(5)
		);
	s_in1(0,5) <= s_out1(1,5);
	s_in2(0,5) <= s_out2(1,6);

		piv_row_6 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,6),
			fetch     => s_fetch(0,6),
			data_in   => s_data_in(0,6),
			data_out  => s_data_out(0,6),
			out1      => s_out1(0,6),
			out2      => s_out2(0,6),
			in1       => s_in1(0,6),
			in2       => s_in2(0,6),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(6)
		);
	s_in1(0,6) <= s_out1(1,6);
	s_in2(0,6) <= s_out2(1,7);

		piv_row_7 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,7),
			fetch     => s_fetch(0,7),
			data_in   => s_data_in(0,7),
			data_out  => s_data_out(0,7),
			out1      => s_out1(0,7),
			out2      => s_out2(0,7),
			in1       => s_in1(0,7),
			in2       => s_in2(0,7),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(7)
		);
	s_in1(0,7) <= s_out1(1,7);
	s_in2(0,7) <= s_out2(1,8);

		piv_row_8 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,8),
			fetch     => s_fetch(0,8),
			data_in   => s_data_in(0,8),
			data_out  => s_data_out(0,8),
			out1      => s_out1(0,8),
			out2      => s_out2(0,8),
			in1       => s_in1(0,8),
			in2       => s_in2(0,8),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(8)
		);
	s_in1(0,8) <= s_out1(1,8);
	s_in2(0,8) <= s_out2(1,9);

		piv_row_9 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,9),
			fetch     => s_fetch(0,9),
			data_in   => s_data_in(0,9),
			data_out  => s_data_out(0,9),
			out1      => s_out1(0,9),
			out2      => s_out2(0,9),
			in1       => s_in1(0,9),
			in2       => s_in2(0,9),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(9)
		);
	s_in1(0,9) <= s_out1(1,9);
	s_in2(0,9) <= s_out2(1,10);

		piv_row_10 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,10),
			fetch     => s_fetch(0,10),
			data_in   => s_data_in(0,10),
			data_out  => s_data_out(0,10),
			out1      => s_out1(0,10),
			out2      => s_out2(0,10),
			in1       => s_in1(0,10),
			in2       => s_in2(0,10),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(10)
		);
	s_in1(0,10) <= s_out1(1,10);
	s_in2(0,10) <= s_out2(1,11);

		piv_row_11 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,11),
			fetch     => s_fetch(0,11),
			data_in   => s_data_in(0,11),
			data_out  => s_data_out(0,11),
			out1      => s_out1(0,11),
			out2      => s_out2(0,11),
			in1       => s_in1(0,11),
			in2       => s_in2(0,11),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(11)
		);
	s_in1(0,11) <= s_out1(1,11);
	s_in2(0,11) <= s_out2(1,12);

		piv_row_12 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,12),
			fetch     => s_fetch(0,12),
			data_in   => s_data_in(0,12),
			data_out  => s_data_out(0,12),
			out1      => s_out1(0,12),
			out2      => s_out2(0,12),
			in1       => s_in1(0,12),
			in2       => s_in2(0,12),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(12)
		);
	s_in1(0,12) <= s_out1(1,12);
	s_in2(0,12) <= s_out2(1,13);

		piv_row_13 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,13),
			fetch     => s_fetch(0,13),
			data_in   => s_data_in(0,13),
			data_out  => s_data_out(0,13),
			out1      => s_out1(0,13),
			out2      => s_out2(0,13),
			in1       => s_in1(0,13),
			in2       => s_in2(0,13),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(13)
		);
	s_in1(0,13) <= s_out1(1,13);
	s_in2(0,13) <= s_out2(1,14);

		piv_row_14 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,14),
			fetch     => s_fetch(0,14),
			data_in   => s_data_in(0,14),
			data_out  => s_data_out(0,14),
			out1      => s_out1(0,14),
			out2      => s_out2(0,14),
			in1       => s_in1(0,14),
			in2       => s_in2(0,14),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(14)
		);
	s_in1(0,14) <= s_out1(1,14);
	s_in2(0,14) <= s_out2(1,15);

		piv_row_15 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,15),
			fetch     => s_fetch(0,15),
			data_in   => s_data_in(0,15),
			data_out  => s_data_out(0,15),
			out1      => s_out1(0,15),
			out2      => s_out2(0,15),
			in1       => s_in1(0,15),
			in2       => s_in2(0,15),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(15)
		);
	s_in1(0,15) <= s_out1(1,15);
	s_in2(0,15) <= s_out2(1,16);

		piv_row_16 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,16),
			fetch     => s_fetch(0,16),
			data_in   => s_data_in(0,16),
			data_out  => s_data_out(0,16),
			out1      => s_out1(0,16),
			out2      => s_out2(0,16),
			in1       => s_in1(0,16),
			in2       => s_in2(0,16),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(16)
		);
	s_in1(0,16) <= s_out1(1,16);
	s_in2(0,16) <= s_out2(1,17);

		piv_row_17 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,17),
			fetch     => s_fetch(0,17),
			data_in   => s_data_in(0,17),
			data_out  => s_data_out(0,17),
			out1      => s_out1(0,17),
			out2      => s_out2(0,17),
			in1       => s_in1(0,17),
			in2       => s_in2(0,17),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(17)
		);
	s_in1(0,17) <= s_out1(1,17);
	s_in2(0,17) <= s_out2(1,18);

		piv_row_18 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,18),
			fetch     => s_fetch(0,18),
			data_in   => s_data_in(0,18),
			data_out  => s_data_out(0,18),
			out1      => s_out1(0,18),
			out2      => s_out2(0,18),
			in1       => s_in1(0,18),
			in2       => s_in2(0,18),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(18)
		);
	s_in1(0,18) <= s_out1(1,18);
	s_in2(0,18) <= s_out2(1,19);

		piv_row_19 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,19),
			fetch     => s_fetch(0,19),
			data_in   => s_data_in(0,19),
			data_out  => s_data_out(0,19),
			out1      => s_out1(0,19),
			out2      => s_out2(0,19),
			in1       => s_in1(0,19),
			in2       => s_in2(0,19),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(19)
		);
	s_in1(0,19) <= s_out1(1,19);
	s_in2(0,19) <= s_out2(1,20);

		piv_row_20 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,20),
			fetch     => s_fetch(0,20),
			data_in   => s_data_in(0,20),
			data_out  => s_data_out(0,20),
			out1      => s_out1(0,20),
			out2      => s_out2(0,20),
			in1       => s_in1(0,20),
			in2       => s_in2(0,20),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(20)
		);
	s_in1(0,20) <= s_out1(1,20);
	s_in2(0,20) <= s_out2(1,21);

		piv_row_21 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,21),
			fetch     => s_fetch(0,21),
			data_in   => s_data_in(0,21),
			data_out  => s_data_out(0,21),
			out1      => s_out1(0,21),
			out2      => s_out2(0,21),
			in1       => s_in1(0,21),
			in2       => s_in2(0,21),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(21)
		);
	s_in1(0,21) <= s_out1(1,21);
	s_in2(0,21) <= s_out2(1,22);

		piv_row_22 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,22),
			fetch     => s_fetch(0,22),
			data_in   => s_data_in(0,22),
			data_out  => s_data_out(0,22),
			out1      => s_out1(0,22),
			out2      => s_out2(0,22),
			in1       => s_in1(0,22),
			in2       => s_in2(0,22),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(22)
		);
	s_in1(0,22) <= s_out1(1,22);
	s_in2(0,22) <= s_out2(1,23);

		piv_row_23 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,23),
			fetch     => s_fetch(0,23),
			data_in   => s_data_in(0,23),
			data_out  => s_data_out(0,23),
			out1      => s_out1(0,23),
			out2      => s_out2(0,23),
			in1       => s_in1(0,23),
			in2       => s_in2(0,23),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(23)
		);
	s_in1(0,23) <= s_out1(1,23);
	s_in2(0,23) <= s_out2(1,24);

		piv_row_24 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,24),
			fetch     => s_fetch(0,24),
			data_in   => s_data_in(0,24),
			data_out  => s_data_out(0,24),
			out1      => s_out1(0,24),
			out2      => s_out2(0,24),
			in1       => s_in1(0,24),
			in2       => s_in2(0,24),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(24)
		);
	s_in1(0,24) <= s_out1(1,24);
	s_in2(0,24) <= s_out2(1,25);

		piv_row_25 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,25),
			fetch     => s_fetch(0,25),
			data_in   => s_data_in(0,25),
			data_out  => s_data_out(0,25),
			out1      => s_out1(0,25),
			out2      => s_out2(0,25),
			in1       => s_in1(0,25),
			in2       => s_in2(0,25),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(25)
		);
	s_in1(0,25) <= s_out1(1,25);
	s_in2(0,25) <= s_out2(1,26);

		piv_row_26 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,26),
			fetch     => s_fetch(0,26),
			data_in   => s_data_in(0,26),
			data_out  => s_data_out(0,26),
			out1      => s_out1(0,26),
			out2      => s_out2(0,26),
			in1       => s_in1(0,26),
			in2       => s_in2(0,26),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(26)
		);
	s_in1(0,26) <= s_out1(1,26);
	s_in2(0,26) <= s_out2(1,27);

		piv_row_27 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,27),
			fetch     => s_fetch(0,27),
			data_in   => s_data_in(0,27),
			data_out  => s_data_out(0,27),
			out1      => s_out1(0,27),
			out2      => s_out2(0,27),
			in1       => s_in1(0,27),
			in2       => s_in2(0,27),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(27)
		);
	s_in1(0,27) <= s_out1(1,27);
	s_in2(0,27) <= s_out2(1,28);

		piv_row_28 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,28),
			fetch     => s_fetch(0,28),
			data_in   => s_data_in(0,28),
			data_out  => s_data_out(0,28),
			out1      => s_out1(0,28),
			out2      => s_out2(0,28),
			in1       => s_in1(0,28),
			in2       => s_in2(0,28),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(28)
		);
	s_in1(0,28) <= s_out1(1,28);
	s_in2(0,28) <= s_out2(1,29);

		piv_row_29 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,29),
			fetch     => s_fetch(0,29),
			data_in   => s_data_in(0,29),
			data_out  => s_data_out(0,29),
			out1      => s_out1(0,29),
			out2      => s_out2(0,29),
			in1       => s_in1(0,29),
			in2       => s_in2(0,29),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(29)
		);
	s_in1(0,29) <= s_out1(1,29);
	s_in2(0,29) <= s_out2(1,30);

		piv_row_30 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,30),
			fetch     => s_fetch(0,30),
			data_in   => s_data_in(0,30),
			data_out  => s_data_out(0,30),
			out1      => s_out1(0,30),
			out2      => s_out2(0,30),
			in1       => s_in1(0,30),
			in2       => s_in2(0,30),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(30)
		);
	s_in1(0,30) <= s_out1(1,30);
	s_in2(0,30) <= s_out2(1,31);

		piv_row_31 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,31),
			fetch     => s_fetch(0,31),
			data_in   => s_data_in(0,31),
			data_out  => s_data_out(0,31),
			out1      => s_out1(0,31),
			out2      => s_out2(0,31),
			in1       => s_in1(0,31),
			in2       => s_in2(0,31),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(31)
		);
	s_in1(0,31) <= s_out1(1,31);
	s_in2(0,31) <= s_out2(1,32);

		piv_row_32 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,32),
			fetch     => s_fetch(0,32),
			data_in   => s_data_in(0,32),
			data_out  => s_data_out(0,32),
			out1      => s_out1(0,32),
			out2      => s_out2(0,32),
			in1       => s_in1(0,32),
			in2       => s_in2(0,32),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(32)
		);
	s_in1(0,32) <= s_out1(1,32);
	s_in2(0,32) <= s_out2(1,33);

		piv_row_33 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,33),
			fetch     => s_fetch(0,33),
			data_in   => s_data_in(0,33),
			data_out  => s_data_out(0,33),
			out1      => s_out1(0,33),
			out2      => s_out2(0,33),
			in1       => s_in1(0,33),
			in2       => s_in2(0,33),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(33)
		);
	s_in1(0,33) <= s_out1(1,33);
	s_in2(0,33) <= s_out2(1,34);

		piv_row_34 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,34),
			fetch     => s_fetch(0,34),
			data_in   => s_data_in(0,34),
			data_out  => s_data_out(0,34),
			out1      => s_out1(0,34),
			out2      => s_out2(0,34),
			in1       => s_in1(0,34),
			in2       => s_in2(0,34),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(34)
		);
	s_in1(0,34) <= s_out1(1,34);
	s_in2(0,34) <= s_out2(1,35);

		piv_row_35 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,35),
			fetch     => s_fetch(0,35),
			data_in   => s_data_in(0,35),
			data_out  => s_data_out(0,35),
			out1      => s_out1(0,35),
			out2      => s_out2(0,35),
			in1       => s_in1(0,35),
			in2       => s_in2(0,35),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(35)
		);
	s_in1(0,35) <= s_out1(1,35);
	s_in2(0,35) <= s_out2(1,36);

		piv_row_36 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,36),
			fetch     => s_fetch(0,36),
			data_in   => s_data_in(0,36),
			data_out  => s_data_out(0,36),
			out1      => s_out1(0,36),
			out2      => s_out2(0,36),
			in1       => s_in1(0,36),
			in2       => s_in2(0,36),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(36)
		);
	s_in1(0,36) <= s_out1(1,36);
	s_in2(0,36) <= s_out2(1,37);

		piv_row_37 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,37),
			fetch     => s_fetch(0,37),
			data_in   => s_data_in(0,37),
			data_out  => s_data_out(0,37),
			out1      => s_out1(0,37),
			out2      => s_out2(0,37),
			in1       => s_in1(0,37),
			in2       => s_in2(0,37),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(37)
		);
	s_in1(0,37) <= s_out1(1,37);
	s_in2(0,37) <= s_out2(1,38);

		piv_row_38 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,38),
			fetch     => s_fetch(0,38),
			data_in   => s_data_in(0,38),
			data_out  => s_data_out(0,38),
			out1      => s_out1(0,38),
			out2      => s_out2(0,38),
			in1       => s_in1(0,38),
			in2       => s_in2(0,38),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(38)
		);
	s_in1(0,38) <= s_out1(1,38);
	s_in2(0,38) <= s_out2(1,39);

		piv_row_39 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,39),
			fetch     => s_fetch(0,39),
			data_in   => s_data_in(0,39),
			data_out  => s_data_out(0,39),
			out1      => s_out1(0,39),
			out2      => s_out2(0,39),
			in1       => s_in1(0,39),
			in2       => s_in2(0,39),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(39)
		);
	s_in1(0,39) <= s_out1(1,39);
	s_in2(0,39) <= s_out2(1,40);

		piv_row_40 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,40),
			fetch     => s_fetch(0,40),
			data_in   => s_data_in(0,40),
			data_out  => s_data_out(0,40),
			out1      => s_out1(0,40),
			out2      => s_out2(0,40),
			in1       => s_in1(0,40),
			in2       => s_in2(0,40),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(40)
		);
	s_in1(0,40) <= s_out1(1,40);
	s_in2(0,40) <= s_out2(1,41);

		piv_row_41 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,41),
			fetch     => s_fetch(0,41),
			data_in   => s_data_in(0,41),
			data_out  => s_data_out(0,41),
			out1      => s_out1(0,41),
			out2      => s_out2(0,41),
			in1       => s_in1(0,41),
			in2       => s_in2(0,41),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(41)
		);
	s_in1(0,41) <= s_out1(1,41);
	s_in2(0,41) <= s_out2(1,42);

		piv_row_42 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,42),
			fetch     => s_fetch(0,42),
			data_in   => s_data_in(0,42),
			data_out  => s_data_out(0,42),
			out1      => s_out1(0,42),
			out2      => s_out2(0,42),
			in1       => s_in1(0,42),
			in2       => s_in2(0,42),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(42)
		);
	s_in1(0,42) <= s_out1(1,42);
	s_in2(0,42) <= s_out2(1,43);

		piv_row_43 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,43),
			fetch     => s_fetch(0,43),
			data_in   => s_data_in(0,43),
			data_out  => s_data_out(0,43),
			out1      => s_out1(0,43),
			out2      => s_out2(0,43),
			in1       => s_in1(0,43),
			in2       => s_in2(0,43),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(43)
		);
	s_in1(0,43) <= s_out1(1,43);
	s_in2(0,43) <= s_out2(1,44);

		piv_row_44 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,44),
			fetch     => s_fetch(0,44),
			data_in   => s_data_in(0,44),
			data_out  => s_data_out(0,44),
			out1      => s_out1(0,44),
			out2      => s_out2(0,44),
			in1       => s_in1(0,44),
			in2       => s_in2(0,44),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(44)
		);
	s_in1(0,44) <= s_out1(1,44);
	s_in2(0,44) <= s_out2(1,45);

		piv_row_45 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,45),
			fetch     => s_fetch(0,45),
			data_in   => s_data_in(0,45),
			data_out  => s_data_out(0,45),
			out1      => s_out1(0,45),
			out2      => s_out2(0,45),
			in1       => s_in1(0,45),
			in2       => s_in2(0,45),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(45)
		);
	s_in1(0,45) <= s_out1(1,45);
	s_in2(0,45) <= s_out2(1,46);

		piv_row_46 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,46),
			fetch     => s_fetch(0,46),
			data_in   => s_data_in(0,46),
			data_out  => s_data_out(0,46),
			out1      => s_out1(0,46),
			out2      => s_out2(0,46),
			in1       => s_in1(0,46),
			in2       => s_in2(0,46),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(46)
		);
	s_in1(0,46) <= s_out1(1,46);
	s_in2(0,46) <= s_out2(1,47);

		piv_row_47 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,47),
			fetch     => s_fetch(0,47),
			data_in   => s_data_in(0,47),
			data_out  => s_data_out(0,47),
			out1      => s_out1(0,47),
			out2      => s_out2(0,47),
			in1       => s_in1(0,47),
			in2       => s_in2(0,47),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(47)
		);
	s_in1(0,47) <= s_out1(1,47);
	s_in2(0,47) <= s_out2(1,48);

		piv_row_48 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,48),
			fetch     => s_fetch(0,48),
			data_in   => s_data_in(0,48),
			data_out  => s_data_out(0,48),
			out1      => s_out1(0,48),
			out2      => s_out2(0,48),
			in1       => s_in1(0,48),
			in2       => s_in2(0,48),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(48)
		);
	s_in1(0,48) <= s_out1(1,48);
	s_in2(0,48) <= s_out2(1,49);

		piv_row_49 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,49),
			fetch     => s_fetch(0,49),
			data_in   => s_data_in(0,49),
			data_out  => s_data_out(0,49),
			out1      => s_out1(0,49),
			out2      => s_out2(0,49),
			in1       => s_in1(0,49),
			in2       => s_in2(0,49),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(49)
		);
	s_in1(0,49) <= s_out1(1,49);
	s_in2(0,49) <= s_out2(1,50);

		piv_row_50 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,50),
			fetch     => s_fetch(0,50),
			data_in   => s_data_in(0,50),
			data_out  => s_data_out(0,50),
			out1      => s_out1(0,50),
			out2      => s_out2(0,50),
			in1       => s_in1(0,50),
			in2       => s_in2(0,50),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(50)
		);
	s_in1(0,50) <= s_out1(1,50);
	s_in2(0,50) <= s_out2(1,51);

		piv_row_51 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,51),
			fetch     => s_fetch(0,51),
			data_in   => s_data_in(0,51),
			data_out  => s_data_out(0,51),
			out1      => s_out1(0,51),
			out2      => s_out2(0,51),
			in1       => s_in1(0,51),
			in2       => s_in2(0,51),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(51)
		);
	s_in1(0,51) <= s_out1(1,51);
	s_in2(0,51) <= s_out2(1,52);

		piv_row_52 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,52),
			fetch     => s_fetch(0,52),
			data_in   => s_data_in(0,52),
			data_out  => s_data_out(0,52),
			out1      => s_out1(0,52),
			out2      => s_out2(0,52),
			in1       => s_in1(0,52),
			in2       => s_in2(0,52),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(52)
		);
	s_in1(0,52) <= s_out1(1,52);
	s_in2(0,52) <= s_out2(1,53);

		piv_row_53 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,53),
			fetch     => s_fetch(0,53),
			data_in   => s_data_in(0,53),
			data_out  => s_data_out(0,53),
			out1      => s_out1(0,53),
			out2      => s_out2(0,53),
			in1       => s_in1(0,53),
			in2       => s_in2(0,53),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(53)
		);
	s_in1(0,53) <= s_out1(1,53);
	s_in2(0,53) <= s_out2(1,54);

		piv_row_54 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,54),
			fetch     => s_fetch(0,54),
			data_in   => s_data_in(0,54),
			data_out  => s_data_out(0,54),
			out1      => s_out1(0,54),
			out2      => s_out2(0,54),
			in1       => s_in1(0,54),
			in2       => s_in2(0,54),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(54)
		);
	s_in1(0,54) <= s_out1(1,54);
	s_in2(0,54) <= s_out2(1,55);

		piv_row_55 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,55),
			fetch     => s_fetch(0,55),
			data_in   => s_data_in(0,55),
			data_out  => s_data_out(0,55),
			out1      => s_out1(0,55),
			out2      => s_out2(0,55),
			in1       => s_in1(0,55),
			in2       => s_in2(0,55),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(55)
		);
	s_in1(0,55) <= s_out1(1,55);
	s_in2(0,55) <= s_out2(1,56);

		piv_row_56 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,56),
			fetch     => s_fetch(0,56),
			data_in   => s_data_in(0,56),
			data_out  => s_data_out(0,56),
			out1      => s_out1(0,56),
			out2      => s_out2(0,56),
			in1       => s_in1(0,56),
			in2       => s_in2(0,56),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(56)
		);
	s_in1(0,56) <= s_out1(1,56);
	s_in2(0,56) <= s_out2(1,57);

		piv_row_57 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,57),
			fetch     => s_fetch(0,57),
			data_in   => s_data_in(0,57),
			data_out  => s_data_out(0,57),
			out1      => s_out1(0,57),
			out2      => s_out2(0,57),
			in1       => s_in1(0,57),
			in2       => s_in2(0,57),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(57)
		);
	s_in1(0,57) <= s_out1(1,57);
	s_in2(0,57) <= s_out2(1,58);

		piv_row_58 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,58),
			fetch     => s_fetch(0,58),
			data_in   => s_data_in(0,58),
			data_out  => s_data_out(0,58),
			out1      => s_out1(0,58),
			out2      => s_out2(0,58),
			in1       => s_in1(0,58),
			in2       => s_in2(0,58),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(58)
		);
	s_in1(0,58) <= s_out1(1,58);
	s_in2(0,58) <= s_out2(1,59);

		piv_row_59 : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,59),
			fetch     => s_fetch(0,59),
			data_in   => s_data_in(0,59),
			data_out  => s_data_out(0,59),
			out1      => s_out1(0,59),
			out2      => s_out2(0,59),
			in1       => s_in1(0,59),
			in2       => s_in2(0,59),
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(59)
		);
	s_in1(0,59) <= s_out1(1,59);
	s_in2(0,59) <= s_out2(1,60);

		piv_row_last : pivotRow_cell port map(
			clk       => clk,
			rst       => rst,
			en        => en,
			load      => s_load(0,60),
			fetch     => s_fetch(0,60),
			data_in   => s_data_in(0,60),
			data_out  => s_data_out(0,60),
			out1      => s_out1(0,COLS-1),
			out2      => s_out2(0,COLS-1),
			in1       => s_in1(0,COLS-1),
			in2       => (others => '0'), -- TODO : Check if cycle is correct
			piv_found => s_piv_found,
			row_data  => s_row_data(0),
			col_data  => s_col_data(COLS-1)
		);
	s_in1(0,60) <= s_out1(1,60);


		--Pivot Cols-----------
		piv_col_1 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,0),
			fetch              => s_fetch(1,0),
			data_in            => s_data_in(1,0),
			data_out           => s_data_out(1,0),
			out1               => s_out1(1,0),
			lock_lower_row_out => s_locks_lower_out(1,0),
			lock_lower_row_in  => s_locks_lower_in(1,0),
			in1                => s_in1(1,0),
			in2                => s_in2(1,0),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1)
		);
	s_in1(1,0)            <= s_out1(2,0);
	s_in2(1,0)            <= s_out2(2,1);
	s_locks_lower_in(1,0) <= s_locks_lower_out(2,0);

		piv_col_2 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,0),
			fetch              => s_fetch(2,0),
			data_in            => s_data_in(2,0),
			data_out           => s_data_out(2,0),
			out1               => s_out1(2,0),
			lock_lower_row_out => s_locks_lower_out(2,0),
			lock_lower_row_in  => s_locks_lower_in(2,0),
			in1                => s_in1(2,0),
			in2                => s_in2(2,0),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2)
		);
	s_in1(2,0)            <= s_out1(3,0);
	s_in2(2,0)            <= s_out2(3,1);
	s_locks_lower_in(2,0) <= s_locks_lower_out(3,0);

		piv_col_3 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,0),
			fetch              => s_fetch(3,0),
			data_in            => s_data_in(3,0),
			data_out           => s_data_out(3,0),
			out1               => s_out1(3,0),
			lock_lower_row_out => s_locks_lower_out(3,0),
			lock_lower_row_in  => s_locks_lower_in(3,0),
			in1                => s_in1(3,0),
			in2                => s_in2(3,0),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3)
		);
	s_in1(3,0)            <= s_out1(4,0);
	s_in2(3,0)            <= s_out2(4,1);
	s_locks_lower_in(3,0) <= s_locks_lower_out(4,0);

		piv_col_4 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,0),
			fetch              => s_fetch(4,0),
			data_in            => s_data_in(4,0),
			data_out           => s_data_out(4,0),
			out1               => s_out1(4,0),
			lock_lower_row_out => s_locks_lower_out(4,0),
			lock_lower_row_in  => s_locks_lower_in(4,0),
			in1                => s_in1(4,0),
			in2                => s_in2(4,0),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4)
		);
	s_in1(4,0)            <= s_out1(5,0);
	s_in2(4,0)            <= s_out2(5,1);
	s_locks_lower_in(4,0) <= s_locks_lower_out(5,0);

		piv_col_5 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,0),
			fetch              => s_fetch(5,0),
			data_in            => s_data_in(5,0),
			data_out           => s_data_out(5,0),
			out1               => s_out1(5,0),
			lock_lower_row_out => s_locks_lower_out(5,0),
			lock_lower_row_in  => s_locks_lower_in(5,0),
			in1                => s_in1(5,0),
			in2                => s_in2(5,0),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5)
		);
	s_in1(5,0)            <= s_out1(6,0);
	s_in2(5,0)            <= s_out2(6,1);
	s_locks_lower_in(5,0) <= s_locks_lower_out(6,0);

		piv_col_6 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,0),
			fetch              => s_fetch(6,0),
			data_in            => s_data_in(6,0),
			data_out           => s_data_out(6,0),
			out1               => s_out1(6,0),
			lock_lower_row_out => s_locks_lower_out(6,0),
			lock_lower_row_in  => s_locks_lower_in(6,0),
			in1                => s_in1(6,0),
			in2                => s_in2(6,0),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6)
		);
	s_in1(6,0)            <= s_out1(7,0);
	s_in2(6,0)            <= s_out2(7,1);
	s_locks_lower_in(6,0) <= s_locks_lower_out(7,0);

		piv_col_7 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,0),
			fetch              => s_fetch(7,0),
			data_in            => s_data_in(7,0),
			data_out           => s_data_out(7,0),
			out1               => s_out1(7,0),
			lock_lower_row_out => s_locks_lower_out(7,0),
			lock_lower_row_in  => s_locks_lower_in(7,0),
			in1                => s_in1(7,0),
			in2                => s_in2(7,0),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7)
		);
	s_in1(7,0)            <= s_out1(8,0);
	s_in2(7,0)            <= s_out2(8,1);
	s_locks_lower_in(7,0) <= s_locks_lower_out(8,0);

		piv_col_8 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,0),
			fetch              => s_fetch(8,0),
			data_in            => s_data_in(8,0),
			data_out           => s_data_out(8,0),
			out1               => s_out1(8,0),
			lock_lower_row_out => s_locks_lower_out(8,0),
			lock_lower_row_in  => s_locks_lower_in(8,0),
			in1                => s_in1(8,0),
			in2                => s_in2(8,0),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8)
		);
	s_in1(8,0)            <= s_out1(9,0);
	s_in2(8,0)            <= s_out2(9,1);
	s_locks_lower_in(8,0) <= s_locks_lower_out(9,0);

		piv_col_9 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,0),
			fetch              => s_fetch(9,0),
			data_in            => s_data_in(9,0),
			data_out           => s_data_out(9,0),
			out1               => s_out1(9,0),
			lock_lower_row_out => s_locks_lower_out(9,0),
			lock_lower_row_in  => s_locks_lower_in(9,0),
			in1                => s_in1(9,0),
			in2                => s_in2(9,0),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9)
		);
	s_in1(9,0)            <= s_out1(10,0);
	s_in2(9,0)            <= s_out2(10,1);
	s_locks_lower_in(9,0) <= s_locks_lower_out(10,0);

		piv_col_10 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,0),
			fetch              => s_fetch(10,0),
			data_in            => s_data_in(10,0),
			data_out           => s_data_out(10,0),
			out1               => s_out1(10,0),
			lock_lower_row_out => s_locks_lower_out(10,0),
			lock_lower_row_in  => s_locks_lower_in(10,0),
			in1                => s_in1(10,0),
			in2                => s_in2(10,0),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10)
		);
	s_in1(10,0)            <= s_out1(11,0);
	s_in2(10,0)            <= s_out2(11,1);
	s_locks_lower_in(10,0) <= s_locks_lower_out(11,0);

		piv_col_11 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,0),
			fetch              => s_fetch(11,0),
			data_in            => s_data_in(11,0),
			data_out           => s_data_out(11,0),
			out1               => s_out1(11,0),
			lock_lower_row_out => s_locks_lower_out(11,0),
			lock_lower_row_in  => s_locks_lower_in(11,0),
			in1                => s_in1(11,0),
			in2                => s_in2(11,0),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11)
		);
	s_in1(11,0)            <= s_out1(12,0);
	s_in2(11,0)            <= s_out2(12,1);
	s_locks_lower_in(11,0) <= s_locks_lower_out(12,0);

		piv_col_12 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,0),
			fetch              => s_fetch(12,0),
			data_in            => s_data_in(12,0),
			data_out           => s_data_out(12,0),
			out1               => s_out1(12,0),
			lock_lower_row_out => s_locks_lower_out(12,0),
			lock_lower_row_in  => s_locks_lower_in(12,0),
			in1                => s_in1(12,0),
			in2                => s_in2(12,0),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12)
		);
	s_in1(12,0)            <= s_out1(13,0);
	s_in2(12,0)            <= s_out2(13,1);
	s_locks_lower_in(12,0) <= s_locks_lower_out(13,0);

		piv_col_13 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,0),
			fetch              => s_fetch(13,0),
			data_in            => s_data_in(13,0),
			data_out           => s_data_out(13,0),
			out1               => s_out1(13,0),
			lock_lower_row_out => s_locks_lower_out(13,0),
			lock_lower_row_in  => s_locks_lower_in(13,0),
			in1                => s_in1(13,0),
			in2                => s_in2(13,0),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13)
		);
	s_in1(13,0)            <= s_out1(14,0);
	s_in2(13,0)            <= s_out2(14,1);
	s_locks_lower_in(13,0) <= s_locks_lower_out(14,0);

		piv_col_14 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,0),
			fetch              => s_fetch(14,0),
			data_in            => s_data_in(14,0),
			data_out           => s_data_out(14,0),
			out1               => s_out1(14,0),
			lock_lower_row_out => s_locks_lower_out(14,0),
			lock_lower_row_in  => s_locks_lower_in(14,0),
			in1                => s_in1(14,0),
			in2                => s_in2(14,0),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14)
		);
	s_in1(14,0)            <= s_out1(15,0);
	s_in2(14,0)            <= s_out2(15,1);
	s_locks_lower_in(14,0) <= s_locks_lower_out(15,0);

		piv_col_15 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,0),
			fetch              => s_fetch(15,0),
			data_in            => s_data_in(15,0),
			data_out           => s_data_out(15,0),
			out1               => s_out1(15,0),
			lock_lower_row_out => s_locks_lower_out(15,0),
			lock_lower_row_in  => s_locks_lower_in(15,0),
			in1                => s_in1(15,0),
			in2                => s_in2(15,0),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15)
		);
	s_in1(15,0)            <= s_out1(16,0);
	s_in2(15,0)            <= s_out2(16,1);
	s_locks_lower_in(15,0) <= s_locks_lower_out(16,0);

		piv_col_16 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,0),
			fetch              => s_fetch(16,0),
			data_in            => s_data_in(16,0),
			data_out           => s_data_out(16,0),
			out1               => s_out1(16,0),
			lock_lower_row_out => s_locks_lower_out(16,0),
			lock_lower_row_in  => s_locks_lower_in(16,0),
			in1                => s_in1(16,0),
			in2                => s_in2(16,0),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16)
		);
	s_in1(16,0)            <= s_out1(17,0);
	s_in2(16,0)            <= s_out2(17,1);
	s_locks_lower_in(16,0) <= s_locks_lower_out(17,0);

		piv_col_17 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,0),
			fetch              => s_fetch(17,0),
			data_in            => s_data_in(17,0),
			data_out           => s_data_out(17,0),
			out1               => s_out1(17,0),
			lock_lower_row_out => s_locks_lower_out(17,0),
			lock_lower_row_in  => s_locks_lower_in(17,0),
			in1                => s_in1(17,0),
			in2                => s_in2(17,0),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17)
		);
	s_in1(17,0)            <= s_out1(18,0);
	s_in2(17,0)            <= s_out2(18,1);
	s_locks_lower_in(17,0) <= s_locks_lower_out(18,0);

		piv_col_18 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,0),
			fetch              => s_fetch(18,0),
			data_in            => s_data_in(18,0),
			data_out           => s_data_out(18,0),
			out1               => s_out1(18,0),
			lock_lower_row_out => s_locks_lower_out(18,0),
			lock_lower_row_in  => s_locks_lower_in(18,0),
			in1                => s_in1(18,0),
			in2                => s_in2(18,0),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18)
		);
	s_in1(18,0)            <= s_out1(19,0);
	s_in2(18,0)            <= s_out2(19,1);
	s_locks_lower_in(18,0) <= s_locks_lower_out(19,0);

		piv_col_19 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,0),
			fetch              => s_fetch(19,0),
			data_in            => s_data_in(19,0),
			data_out           => s_data_out(19,0),
			out1               => s_out1(19,0),
			lock_lower_row_out => s_locks_lower_out(19,0),
			lock_lower_row_in  => s_locks_lower_in(19,0),
			in1                => s_in1(19,0),
			in2                => s_in2(19,0),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19)
		);
	s_in1(19,0)            <= s_out1(20,0);
	s_in2(19,0)            <= s_out2(20,1);
	s_locks_lower_in(19,0) <= s_locks_lower_out(20,0);

		piv_col_20 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,0),
			fetch              => s_fetch(20,0),
			data_in            => s_data_in(20,0),
			data_out           => s_data_out(20,0),
			out1               => s_out1(20,0),
			lock_lower_row_out => s_locks_lower_out(20,0),
			lock_lower_row_in  => s_locks_lower_in(20,0),
			in1                => s_in1(20,0),
			in2                => s_in2(20,0),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20)
		);
	s_in1(20,0)            <= s_out1(21,0);
	s_in2(20,0)            <= s_out2(21,1);
	s_locks_lower_in(20,0) <= s_locks_lower_out(21,0);

		piv_col_21 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,0),
			fetch              => s_fetch(21,0),
			data_in            => s_data_in(21,0),
			data_out           => s_data_out(21,0),
			out1               => s_out1(21,0),
			lock_lower_row_out => s_locks_lower_out(21,0),
			lock_lower_row_in  => s_locks_lower_in(21,0),
			in1                => s_in1(21,0),
			in2                => s_in2(21,0),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21)
		);
	s_in1(21,0)            <= s_out1(22,0);
	s_in2(21,0)            <= s_out2(22,1);
	s_locks_lower_in(21,0) <= s_locks_lower_out(22,0);

		piv_col_22 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,0),
			fetch              => s_fetch(22,0),
			data_in            => s_data_in(22,0),
			data_out           => s_data_out(22,0),
			out1               => s_out1(22,0),
			lock_lower_row_out => s_locks_lower_out(22,0),
			lock_lower_row_in  => s_locks_lower_in(22,0),
			in1                => s_in1(22,0),
			in2                => s_in2(22,0),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22)
		);
	s_in1(22,0)            <= s_out1(23,0);
	s_in2(22,0)            <= s_out2(23,1);
	s_locks_lower_in(22,0) <= s_locks_lower_out(23,0);

		piv_col_23 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,0),
			fetch              => s_fetch(23,0),
			data_in            => s_data_in(23,0),
			data_out           => s_data_out(23,0),
			out1               => s_out1(23,0),
			lock_lower_row_out => s_locks_lower_out(23,0),
			lock_lower_row_in  => s_locks_lower_in(23,0),
			in1                => s_in1(23,0),
			in2                => s_in2(23,0),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23)
		);
	s_in1(23,0)            <= s_out1(24,0);
	s_in2(23,0)            <= s_out2(24,1);
	s_locks_lower_in(23,0) <= s_locks_lower_out(24,0);

		piv_col_24 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,0),
			fetch              => s_fetch(24,0),
			data_in            => s_data_in(24,0),
			data_out           => s_data_out(24,0),
			out1               => s_out1(24,0),
			lock_lower_row_out => s_locks_lower_out(24,0),
			lock_lower_row_in  => s_locks_lower_in(24,0),
			in1                => s_in1(24,0),
			in2                => s_in2(24,0),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24)
		);
	s_in1(24,0)            <= s_out1(25,0);
	s_in2(24,0)            <= s_out2(25,1);
	s_locks_lower_in(24,0) <= s_locks_lower_out(25,0);

		piv_col_25 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,0),
			fetch              => s_fetch(25,0),
			data_in            => s_data_in(25,0),
			data_out           => s_data_out(25,0),
			out1               => s_out1(25,0),
			lock_lower_row_out => s_locks_lower_out(25,0),
			lock_lower_row_in  => s_locks_lower_in(25,0),
			in1                => s_in1(25,0),
			in2                => s_in2(25,0),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25)
		);
	s_in1(25,0)            <= s_out1(26,0);
	s_in2(25,0)            <= s_out2(26,1);
	s_locks_lower_in(25,0) <= s_locks_lower_out(26,0);

		piv_col_26 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,0),
			fetch              => s_fetch(26,0),
			data_in            => s_data_in(26,0),
			data_out           => s_data_out(26,0),
			out1               => s_out1(26,0),
			lock_lower_row_out => s_locks_lower_out(26,0),
			lock_lower_row_in  => s_locks_lower_in(26,0),
			in1                => s_in1(26,0),
			in2                => s_in2(26,0),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26)
		);
	s_in1(26,0)            <= s_out1(27,0);
	s_in2(26,0)            <= s_out2(27,1);
	s_locks_lower_in(26,0) <= s_locks_lower_out(27,0);

		piv_col_27 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,0),
			fetch              => s_fetch(27,0),
			data_in            => s_data_in(27,0),
			data_out           => s_data_out(27,0),
			out1               => s_out1(27,0),
			lock_lower_row_out => s_locks_lower_out(27,0),
			lock_lower_row_in  => s_locks_lower_in(27,0),
			in1                => s_in1(27,0),
			in2                => s_in2(27,0),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27)
		);
	s_in1(27,0)            <= s_out1(28,0);
	s_in2(27,0)            <= s_out2(28,1);
	s_locks_lower_in(27,0) <= s_locks_lower_out(28,0);

		piv_col_28 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,0),
			fetch              => s_fetch(28,0),
			data_in            => s_data_in(28,0),
			data_out           => s_data_out(28,0),
			out1               => s_out1(28,0),
			lock_lower_row_out => s_locks_lower_out(28,0),
			lock_lower_row_in  => s_locks_lower_in(28,0),
			in1                => s_in1(28,0),
			in2                => s_in2(28,0),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28)
		);
	s_in1(28,0)            <= s_out1(29,0);
	s_in2(28,0)            <= s_out2(29,1);
	s_locks_lower_in(28,0) <= s_locks_lower_out(29,0);

		piv_col_29 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,0),
			fetch              => s_fetch(29,0),
			data_in            => s_data_in(29,0),
			data_out           => s_data_out(29,0),
			out1               => s_out1(29,0),
			lock_lower_row_out => s_locks_lower_out(29,0),
			lock_lower_row_in  => s_locks_lower_in(29,0),
			in1                => s_in1(29,0),
			in2                => s_in2(29,0),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29)
		);
	s_in1(29,0)            <= s_out1(30,0);
	s_in2(29,0)            <= s_out2(30,1);
	s_locks_lower_in(29,0) <= s_locks_lower_out(30,0);

		piv_col_30 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,0),
			fetch              => s_fetch(30,0),
			data_in            => s_data_in(30,0),
			data_out           => s_data_out(30,0),
			out1               => s_out1(30,0),
			lock_lower_row_out => s_locks_lower_out(30,0),
			lock_lower_row_in  => s_locks_lower_in(30,0),
			in1                => s_in1(30,0),
			in2                => s_in2(30,0),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30)
		);
	s_in1(30,0)            <= s_out1(31,0);
	s_in2(30,0)            <= s_out2(31,1);
	s_locks_lower_in(30,0) <= s_locks_lower_out(31,0);

		piv_col_31 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,0),
			fetch              => s_fetch(31,0),
			data_in            => s_data_in(31,0),
			data_out           => s_data_out(31,0),
			out1               => s_out1(31,0),
			lock_lower_row_out => s_locks_lower_out(31,0),
			lock_lower_row_in  => s_locks_lower_in(31,0),
			in1                => s_in1(31,0),
			in2                => s_in2(31,0),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31)
		);
	s_in1(31,0)            <= s_out1(32,0);
	s_in2(31,0)            <= s_out2(32,1);
	s_locks_lower_in(31,0) <= s_locks_lower_out(32,0);

		piv_col_32 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,0),
			fetch              => s_fetch(32,0),
			data_in            => s_data_in(32,0),
			data_out           => s_data_out(32,0),
			out1               => s_out1(32,0),
			lock_lower_row_out => s_locks_lower_out(32,0),
			lock_lower_row_in  => s_locks_lower_in(32,0),
			in1                => s_in1(32,0),
			in2                => s_in2(32,0),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32)
		);
	s_in1(32,0)            <= s_out1(33,0);
	s_in2(32,0)            <= s_out2(33,1);
	s_locks_lower_in(32,0) <= s_locks_lower_out(33,0);

		piv_col_33 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,0),
			fetch              => s_fetch(33,0),
			data_in            => s_data_in(33,0),
			data_out           => s_data_out(33,0),
			out1               => s_out1(33,0),
			lock_lower_row_out => s_locks_lower_out(33,0),
			lock_lower_row_in  => s_locks_lower_in(33,0),
			in1                => s_in1(33,0),
			in2                => s_in2(33,0),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33)
		);
	s_in1(33,0)            <= s_out1(34,0);
	s_in2(33,0)            <= s_out2(34,1);
	s_locks_lower_in(33,0) <= s_locks_lower_out(34,0);

		piv_col_34 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,0),
			fetch              => s_fetch(34,0),
			data_in            => s_data_in(34,0),
			data_out           => s_data_out(34,0),
			out1               => s_out1(34,0),
			lock_lower_row_out => s_locks_lower_out(34,0),
			lock_lower_row_in  => s_locks_lower_in(34,0),
			in1                => s_in1(34,0),
			in2                => s_in2(34,0),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34)
		);
	s_in1(34,0)            <= s_out1(35,0);
	s_in2(34,0)            <= s_out2(35,1);
	s_locks_lower_in(34,0) <= s_locks_lower_out(35,0);

		piv_col_35 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,0),
			fetch              => s_fetch(35,0),
			data_in            => s_data_in(35,0),
			data_out           => s_data_out(35,0),
			out1               => s_out1(35,0),
			lock_lower_row_out => s_locks_lower_out(35,0),
			lock_lower_row_in  => s_locks_lower_in(35,0),
			in1                => s_in1(35,0),
			in2                => s_in2(35,0),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35)
		);
	s_in1(35,0)            <= s_out1(36,0);
	s_in2(35,0)            <= s_out2(36,1);
	s_locks_lower_in(35,0) <= s_locks_lower_out(36,0);

		piv_col_36 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,0),
			fetch              => s_fetch(36,0),
			data_in            => s_data_in(36,0),
			data_out           => s_data_out(36,0),
			out1               => s_out1(36,0),
			lock_lower_row_out => s_locks_lower_out(36,0),
			lock_lower_row_in  => s_locks_lower_in(36,0),
			in1                => s_in1(36,0),
			in2                => s_in2(36,0),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36)
		);
	s_in1(36,0)            <= s_out1(37,0);
	s_in2(36,0)            <= s_out2(37,1);
	s_locks_lower_in(36,0) <= s_locks_lower_out(37,0);

		piv_col_37 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,0),
			fetch              => s_fetch(37,0),
			data_in            => s_data_in(37,0),
			data_out           => s_data_out(37,0),
			out1               => s_out1(37,0),
			lock_lower_row_out => s_locks_lower_out(37,0),
			lock_lower_row_in  => s_locks_lower_in(37,0),
			in1                => s_in1(37,0),
			in2                => s_in2(37,0),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37)
		);
	s_in1(37,0)            <= s_out1(38,0);
	s_in2(37,0)            <= s_out2(38,1);
	s_locks_lower_in(37,0) <= s_locks_lower_out(38,0);

		piv_col_38 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,0),
			fetch              => s_fetch(38,0),
			data_in            => s_data_in(38,0),
			data_out           => s_data_out(38,0),
			out1               => s_out1(38,0),
			lock_lower_row_out => s_locks_lower_out(38,0),
			lock_lower_row_in  => s_locks_lower_in(38,0),
			in1                => s_in1(38,0),
			in2                => s_in2(38,0),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38)
		);
	s_in1(38,0)            <= s_out1(39,0);
	s_in2(38,0)            <= s_out2(39,1);
	s_locks_lower_in(38,0) <= s_locks_lower_out(39,0);

		piv_col_39 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,0),
			fetch              => s_fetch(39,0),
			data_in            => s_data_in(39,0),
			data_out           => s_data_out(39,0),
			out1               => s_out1(39,0),
			lock_lower_row_out => s_locks_lower_out(39,0),
			lock_lower_row_in  => s_locks_lower_in(39,0),
			in1                => s_in1(39,0),
			in2                => s_in2(39,0),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39)
		);
	s_in1(39,0)            <= s_out1(40,0);
	s_in2(39,0)            <= s_out2(40,1);
	s_locks_lower_in(39,0) <= s_locks_lower_out(40,0);

		piv_col_40 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,0),
			fetch              => s_fetch(40,0),
			data_in            => s_data_in(40,0),
			data_out           => s_data_out(40,0),
			out1               => s_out1(40,0),
			lock_lower_row_out => s_locks_lower_out(40,0),
			lock_lower_row_in  => s_locks_lower_in(40,0),
			in1                => s_in1(40,0),
			in2                => s_in2(40,0),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40)
		);
	s_in1(40,0)            <= s_out1(41,0);
	s_in2(40,0)            <= s_out2(41,1);
	s_locks_lower_in(40,0) <= s_locks_lower_out(41,0);

		piv_col_41 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,0),
			fetch              => s_fetch(41,0),
			data_in            => s_data_in(41,0),
			data_out           => s_data_out(41,0),
			out1               => s_out1(41,0),
			lock_lower_row_out => s_locks_lower_out(41,0),
			lock_lower_row_in  => s_locks_lower_in(41,0),
			in1                => s_in1(41,0),
			in2                => s_in2(41,0),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41)
		);
	s_in1(41,0)            <= s_out1(42,0);
	s_in2(41,0)            <= s_out2(42,1);
	s_locks_lower_in(41,0) <= s_locks_lower_out(42,0);

		piv_col_42 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,0),
			fetch              => s_fetch(42,0),
			data_in            => s_data_in(42,0),
			data_out           => s_data_out(42,0),
			out1               => s_out1(42,0),
			lock_lower_row_out => s_locks_lower_out(42,0),
			lock_lower_row_in  => s_locks_lower_in(42,0),
			in1                => s_in1(42,0),
			in2                => s_in2(42,0),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42)
		);
	s_in1(42,0)            <= s_out1(43,0);
	s_in2(42,0)            <= s_out2(43,1);
	s_locks_lower_in(42,0) <= s_locks_lower_out(43,0);

		piv_col_43 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,0),
			fetch              => s_fetch(43,0),
			data_in            => s_data_in(43,0),
			data_out           => s_data_out(43,0),
			out1               => s_out1(43,0),
			lock_lower_row_out => s_locks_lower_out(43,0),
			lock_lower_row_in  => s_locks_lower_in(43,0),
			in1                => s_in1(43,0),
			in2                => s_in2(43,0),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43)
		);
	s_in1(43,0)            <= s_out1(44,0);
	s_in2(43,0)            <= s_out2(44,1);
	s_locks_lower_in(43,0) <= s_locks_lower_out(44,0);

		piv_col_44 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,0),
			fetch              => s_fetch(44,0),
			data_in            => s_data_in(44,0),
			data_out           => s_data_out(44,0),
			out1               => s_out1(44,0),
			lock_lower_row_out => s_locks_lower_out(44,0),
			lock_lower_row_in  => s_locks_lower_in(44,0),
			in1                => s_in1(44,0),
			in2                => s_in2(44,0),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44)
		);
	s_in1(44,0)            <= s_out1(45,0);
	s_in2(44,0)            <= s_out2(45,1);
	s_locks_lower_in(44,0) <= s_locks_lower_out(45,0);

		piv_col_45 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,0),
			fetch              => s_fetch(45,0),
			data_in            => s_data_in(45,0),
			data_out           => s_data_out(45,0),
			out1               => s_out1(45,0),
			lock_lower_row_out => s_locks_lower_out(45,0),
			lock_lower_row_in  => s_locks_lower_in(45,0),
			in1                => s_in1(45,0),
			in2                => s_in2(45,0),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45)
		);
	s_in1(45,0)            <= s_out1(46,0);
	s_in2(45,0)            <= s_out2(46,1);
	s_locks_lower_in(45,0) <= s_locks_lower_out(46,0);

		piv_col_46 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,0),
			fetch              => s_fetch(46,0),
			data_in            => s_data_in(46,0),
			data_out           => s_data_out(46,0),
			out1               => s_out1(46,0),
			lock_lower_row_out => s_locks_lower_out(46,0),
			lock_lower_row_in  => s_locks_lower_in(46,0),
			in1                => s_in1(46,0),
			in2                => s_in2(46,0),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46)
		);
	s_in1(46,0)            <= s_out1(47,0);
	s_in2(46,0)            <= s_out2(47,1);
	s_locks_lower_in(46,0) <= s_locks_lower_out(47,0);

		piv_col_47 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,0),
			fetch              => s_fetch(47,0),
			data_in            => s_data_in(47,0),
			data_out           => s_data_out(47,0),
			out1               => s_out1(47,0),
			lock_lower_row_out => s_locks_lower_out(47,0),
			lock_lower_row_in  => s_locks_lower_in(47,0),
			in1                => s_in1(47,0),
			in2                => s_in2(47,0),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47)
		);
	s_in1(47,0)            <= s_out1(48,0);
	s_in2(47,0)            <= s_out2(48,1);
	s_locks_lower_in(47,0) <= s_locks_lower_out(48,0);

		piv_col_48 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,0),
			fetch              => s_fetch(48,0),
			data_in            => s_data_in(48,0),
			data_out           => s_data_out(48,0),
			out1               => s_out1(48,0),
			lock_lower_row_out => s_locks_lower_out(48,0),
			lock_lower_row_in  => s_locks_lower_in(48,0),
			in1                => s_in1(48,0),
			in2                => s_in2(48,0),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48)
		);
	s_in1(48,0)            <= s_out1(49,0);
	s_in2(48,0)            <= s_out2(49,1);
	s_locks_lower_in(48,0) <= s_locks_lower_out(49,0);

		piv_col_49 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,0),
			fetch              => s_fetch(49,0),
			data_in            => s_data_in(49,0),
			data_out           => s_data_out(49,0),
			out1               => s_out1(49,0),
			lock_lower_row_out => s_locks_lower_out(49,0),
			lock_lower_row_in  => s_locks_lower_in(49,0),
			in1                => s_in1(49,0),
			in2                => s_in2(49,0),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49)
		);
	s_in1(49,0)            <= s_out1(50,0);
	s_in2(49,0)            <= s_out2(50,1);
	s_locks_lower_in(49,0) <= s_locks_lower_out(50,0);

		piv_col_50 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,0),
			fetch              => s_fetch(50,0),
			data_in            => s_data_in(50,0),
			data_out           => s_data_out(50,0),
			out1               => s_out1(50,0),
			lock_lower_row_out => s_locks_lower_out(50,0),
			lock_lower_row_in  => s_locks_lower_in(50,0),
			in1                => s_in1(50,0),
			in2                => s_in2(50,0),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50)
		);
	s_in1(50,0)            <= s_out1(51,0);
	s_in2(50,0)            <= s_out2(51,1);
	s_locks_lower_in(50,0) <= s_locks_lower_out(51,0);

		piv_col_51 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,0),
			fetch              => s_fetch(51,0),
			data_in            => s_data_in(51,0),
			data_out           => s_data_out(51,0),
			out1               => s_out1(51,0),
			lock_lower_row_out => s_locks_lower_out(51,0),
			lock_lower_row_in  => s_locks_lower_in(51,0),
			in1                => s_in1(51,0),
			in2                => s_in2(51,0),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51)
		);
	s_in1(51,0)            <= s_out1(52,0);
	s_in2(51,0)            <= s_out2(52,1);
	s_locks_lower_in(51,0) <= s_locks_lower_out(52,0);

		piv_col_52 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,0),
			fetch              => s_fetch(52,0),
			data_in            => s_data_in(52,0),
			data_out           => s_data_out(52,0),
			out1               => s_out1(52,0),
			lock_lower_row_out => s_locks_lower_out(52,0),
			lock_lower_row_in  => s_locks_lower_in(52,0),
			in1                => s_in1(52,0),
			in2                => s_in2(52,0),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52)
		);
	s_in1(52,0)            <= s_out1(53,0);
	s_in2(52,0)            <= s_out2(53,1);
	s_locks_lower_in(52,0) <= s_locks_lower_out(53,0);

		piv_col_53 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,0),
			fetch              => s_fetch(53,0),
			data_in            => s_data_in(53,0),
			data_out           => s_data_out(53,0),
			out1               => s_out1(53,0),
			lock_lower_row_out => s_locks_lower_out(53,0),
			lock_lower_row_in  => s_locks_lower_in(53,0),
			in1                => s_in1(53,0),
			in2                => s_in2(53,0),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53)
		);
	s_in1(53,0)            <= s_out1(54,0);
	s_in2(53,0)            <= s_out2(54,1);
	s_locks_lower_in(53,0) <= s_locks_lower_out(54,0);

		piv_col_54 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,0),
			fetch              => s_fetch(54,0),
			data_in            => s_data_in(54,0),
			data_out           => s_data_out(54,0),
			out1               => s_out1(54,0),
			lock_lower_row_out => s_locks_lower_out(54,0),
			lock_lower_row_in  => s_locks_lower_in(54,0),
			in1                => s_in1(54,0),
			in2                => s_in2(54,0),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54)
		);
	s_in1(54,0)            <= s_out1(55,0);
	s_in2(54,0)            <= s_out2(55,1);
	s_locks_lower_in(54,0) <= s_locks_lower_out(55,0);

		piv_col_55 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,0),
			fetch              => s_fetch(55,0),
			data_in            => s_data_in(55,0),
			data_out           => s_data_out(55,0),
			out1               => s_out1(55,0),
			lock_lower_row_out => s_locks_lower_out(55,0),
			lock_lower_row_in  => s_locks_lower_in(55,0),
			in1                => s_in1(55,0),
			in2                => s_in2(55,0),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55)
		);
	s_in1(55,0)            <= s_out1(56,0);
	s_in2(55,0)            <= s_out2(56,1);
	s_locks_lower_in(55,0) <= s_locks_lower_out(56,0);

		piv_col_56 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,0),
			fetch              => s_fetch(56,0),
			data_in            => s_data_in(56,0),
			data_out           => s_data_out(56,0),
			out1               => s_out1(56,0),
			lock_lower_row_out => s_locks_lower_out(56,0),
			lock_lower_row_in  => s_locks_lower_in(56,0),
			in1                => s_in1(56,0),
			in2                => s_in2(56,0),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56)
		);
	s_in1(56,0)            <= s_out1(57,0);
	s_in2(56,0)            <= s_out2(57,1);
	s_locks_lower_in(56,0) <= s_locks_lower_out(57,0);

		piv_col_57 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,0),
			fetch              => s_fetch(57,0),
			data_in            => s_data_in(57,0),
			data_out           => s_data_out(57,0),
			out1               => s_out1(57,0),
			lock_lower_row_out => s_locks_lower_out(57,0),
			lock_lower_row_in  => s_locks_lower_in(57,0),
			in1                => s_in1(57,0),
			in2                => s_in2(57,0),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57)
		);
	s_in1(57,0)            <= s_out1(58,0);
	s_in2(57,0)            <= s_out2(58,1);
	s_locks_lower_in(57,0) <= s_locks_lower_out(58,0);

		piv_col_58 : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,0),
			fetch              => s_fetch(58,0),
			data_in            => s_data_in(58,0),
			data_out           => s_data_out(58,0),
			out1               => s_out1(58,0),
			lock_lower_row_out => s_locks_lower_out(58,0),
			lock_lower_row_in  => s_locks_lower_in(58,0),
			in1                => s_in1(58,0),
			in2                => s_in2(58,0),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58)
		);
	s_in1(58,0)            <= s_out1(59,0);
	s_in2(58,0)            <= s_out2(59,1);
	s_locks_lower_in(58,0) <= s_locks_lower_out(59,0);

		last_piv_col : pivotCol_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,0),
			fetch              => s_fetch(59,0),
			data_in            => s_data_in(59,0),
			data_out           => s_data_out(59,0),
			out1               => s_out1(59,0),
			lock_lower_row_out => s_locks_lower_out(59,0),
			lock_lower_row_in  => '0',
			in1                => (others => '0'),
			in2                => s_in2(59,0),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59)
		);
	s_in2(59,0) <= s_out2(0,1);


		--Basic Cells----------
		normal_cell_1_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,1),
			fetch              => s_fetch(1,1),
			data_in            => s_data_in(1,1),
			data_out           => s_data_out(1,1),
			out1               => s_out1(1,1),
			out2               => s_out2(1,1),
			lock_lower_row_out => s_locks_lower_out(1,1),
			lock_lower_row_in  => s_locks_lower_in(1,1),
			in1                => s_in1(1,1),
			in2                => s_in2(1,1),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(1)
		);
	s_in1(1,1)            <= s_out1(2,1);
	s_in2(1,1)            <= s_out2(2,2);
	s_locks_lower_in(1,1) <= s_locks_lower_out(2,1);

		normal_cell_1_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,2),
			fetch              => s_fetch(1,2),
			data_in            => s_data_in(1,2),
			data_out           => s_data_out(1,2),
			out1               => s_out1(1,2),
			out2               => s_out2(1,2),
			lock_lower_row_out => s_locks_lower_out(1,2),
			lock_lower_row_in  => s_locks_lower_in(1,2),
			in1                => s_in1(1,2),
			in2                => s_in2(1,2),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(2)
		);
	s_in1(1,2)            <= s_out1(2,2);
	s_in2(1,2)            <= s_out2(2,3);
	s_locks_lower_in(1,2) <= s_locks_lower_out(2,2);

		normal_cell_1_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,3),
			fetch              => s_fetch(1,3),
			data_in            => s_data_in(1,3),
			data_out           => s_data_out(1,3),
			out1               => s_out1(1,3),
			out2               => s_out2(1,3),
			lock_lower_row_out => s_locks_lower_out(1,3),
			lock_lower_row_in  => s_locks_lower_in(1,3),
			in1                => s_in1(1,3),
			in2                => s_in2(1,3),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(3)
		);
	s_in1(1,3)            <= s_out1(2,3);
	s_in2(1,3)            <= s_out2(2,4);
	s_locks_lower_in(1,3) <= s_locks_lower_out(2,3);

		normal_cell_1_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,4),
			fetch              => s_fetch(1,4),
			data_in            => s_data_in(1,4),
			data_out           => s_data_out(1,4),
			out1               => s_out1(1,4),
			out2               => s_out2(1,4),
			lock_lower_row_out => s_locks_lower_out(1,4),
			lock_lower_row_in  => s_locks_lower_in(1,4),
			in1                => s_in1(1,4),
			in2                => s_in2(1,4),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(4)
		);
	s_in1(1,4)            <= s_out1(2,4);
	s_in2(1,4)            <= s_out2(2,5);
	s_locks_lower_in(1,4) <= s_locks_lower_out(2,4);

		normal_cell_1_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,5),
			fetch              => s_fetch(1,5),
			data_in            => s_data_in(1,5),
			data_out           => s_data_out(1,5),
			out1               => s_out1(1,5),
			out2               => s_out2(1,5),
			lock_lower_row_out => s_locks_lower_out(1,5),
			lock_lower_row_in  => s_locks_lower_in(1,5),
			in1                => s_in1(1,5),
			in2                => s_in2(1,5),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(5)
		);
	s_in1(1,5)            <= s_out1(2,5);
	s_in2(1,5)            <= s_out2(2,6);
	s_locks_lower_in(1,5) <= s_locks_lower_out(2,5);

		normal_cell_1_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,6),
			fetch              => s_fetch(1,6),
			data_in            => s_data_in(1,6),
			data_out           => s_data_out(1,6),
			out1               => s_out1(1,6),
			out2               => s_out2(1,6),
			lock_lower_row_out => s_locks_lower_out(1,6),
			lock_lower_row_in  => s_locks_lower_in(1,6),
			in1                => s_in1(1,6),
			in2                => s_in2(1,6),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(6)
		);
	s_in1(1,6)            <= s_out1(2,6);
	s_in2(1,6)            <= s_out2(2,7);
	s_locks_lower_in(1,6) <= s_locks_lower_out(2,6);

		normal_cell_1_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,7),
			fetch              => s_fetch(1,7),
			data_in            => s_data_in(1,7),
			data_out           => s_data_out(1,7),
			out1               => s_out1(1,7),
			out2               => s_out2(1,7),
			lock_lower_row_out => s_locks_lower_out(1,7),
			lock_lower_row_in  => s_locks_lower_in(1,7),
			in1                => s_in1(1,7),
			in2                => s_in2(1,7),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(7)
		);
	s_in1(1,7)            <= s_out1(2,7);
	s_in2(1,7)            <= s_out2(2,8);
	s_locks_lower_in(1,7) <= s_locks_lower_out(2,7);

		normal_cell_1_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,8),
			fetch              => s_fetch(1,8),
			data_in            => s_data_in(1,8),
			data_out           => s_data_out(1,8),
			out1               => s_out1(1,8),
			out2               => s_out2(1,8),
			lock_lower_row_out => s_locks_lower_out(1,8),
			lock_lower_row_in  => s_locks_lower_in(1,8),
			in1                => s_in1(1,8),
			in2                => s_in2(1,8),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(8)
		);
	s_in1(1,8)            <= s_out1(2,8);
	s_in2(1,8)            <= s_out2(2,9);
	s_locks_lower_in(1,8) <= s_locks_lower_out(2,8);

		normal_cell_1_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,9),
			fetch              => s_fetch(1,9),
			data_in            => s_data_in(1,9),
			data_out           => s_data_out(1,9),
			out1               => s_out1(1,9),
			out2               => s_out2(1,9),
			lock_lower_row_out => s_locks_lower_out(1,9),
			lock_lower_row_in  => s_locks_lower_in(1,9),
			in1                => s_in1(1,9),
			in2                => s_in2(1,9),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(9)
		);
	s_in1(1,9)            <= s_out1(2,9);
	s_in2(1,9)            <= s_out2(2,10);
	s_locks_lower_in(1,9) <= s_locks_lower_out(2,9);

		normal_cell_1_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,10),
			fetch              => s_fetch(1,10),
			data_in            => s_data_in(1,10),
			data_out           => s_data_out(1,10),
			out1               => s_out1(1,10),
			out2               => s_out2(1,10),
			lock_lower_row_out => s_locks_lower_out(1,10),
			lock_lower_row_in  => s_locks_lower_in(1,10),
			in1                => s_in1(1,10),
			in2                => s_in2(1,10),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(10)
		);
	s_in1(1,10)            <= s_out1(2,10);
	s_in2(1,10)            <= s_out2(2,11);
	s_locks_lower_in(1,10) <= s_locks_lower_out(2,10);

		normal_cell_1_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,11),
			fetch              => s_fetch(1,11),
			data_in            => s_data_in(1,11),
			data_out           => s_data_out(1,11),
			out1               => s_out1(1,11),
			out2               => s_out2(1,11),
			lock_lower_row_out => s_locks_lower_out(1,11),
			lock_lower_row_in  => s_locks_lower_in(1,11),
			in1                => s_in1(1,11),
			in2                => s_in2(1,11),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(11)
		);
	s_in1(1,11)            <= s_out1(2,11);
	s_in2(1,11)            <= s_out2(2,12);
	s_locks_lower_in(1,11) <= s_locks_lower_out(2,11);

		normal_cell_1_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,12),
			fetch              => s_fetch(1,12),
			data_in            => s_data_in(1,12),
			data_out           => s_data_out(1,12),
			out1               => s_out1(1,12),
			out2               => s_out2(1,12),
			lock_lower_row_out => s_locks_lower_out(1,12),
			lock_lower_row_in  => s_locks_lower_in(1,12),
			in1                => s_in1(1,12),
			in2                => s_in2(1,12),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(12)
		);
	s_in1(1,12)            <= s_out1(2,12);
	s_in2(1,12)            <= s_out2(2,13);
	s_locks_lower_in(1,12) <= s_locks_lower_out(2,12);

		normal_cell_1_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,13),
			fetch              => s_fetch(1,13),
			data_in            => s_data_in(1,13),
			data_out           => s_data_out(1,13),
			out1               => s_out1(1,13),
			out2               => s_out2(1,13),
			lock_lower_row_out => s_locks_lower_out(1,13),
			lock_lower_row_in  => s_locks_lower_in(1,13),
			in1                => s_in1(1,13),
			in2                => s_in2(1,13),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(13)
		);
	s_in1(1,13)            <= s_out1(2,13);
	s_in2(1,13)            <= s_out2(2,14);
	s_locks_lower_in(1,13) <= s_locks_lower_out(2,13);

		normal_cell_1_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,14),
			fetch              => s_fetch(1,14),
			data_in            => s_data_in(1,14),
			data_out           => s_data_out(1,14),
			out1               => s_out1(1,14),
			out2               => s_out2(1,14),
			lock_lower_row_out => s_locks_lower_out(1,14),
			lock_lower_row_in  => s_locks_lower_in(1,14),
			in1                => s_in1(1,14),
			in2                => s_in2(1,14),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(14)
		);
	s_in1(1,14)            <= s_out1(2,14);
	s_in2(1,14)            <= s_out2(2,15);
	s_locks_lower_in(1,14) <= s_locks_lower_out(2,14);

		normal_cell_1_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,15),
			fetch              => s_fetch(1,15),
			data_in            => s_data_in(1,15),
			data_out           => s_data_out(1,15),
			out1               => s_out1(1,15),
			out2               => s_out2(1,15),
			lock_lower_row_out => s_locks_lower_out(1,15),
			lock_lower_row_in  => s_locks_lower_in(1,15),
			in1                => s_in1(1,15),
			in2                => s_in2(1,15),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(15)
		);
	s_in1(1,15)            <= s_out1(2,15);
	s_in2(1,15)            <= s_out2(2,16);
	s_locks_lower_in(1,15) <= s_locks_lower_out(2,15);

		normal_cell_1_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,16),
			fetch              => s_fetch(1,16),
			data_in            => s_data_in(1,16),
			data_out           => s_data_out(1,16),
			out1               => s_out1(1,16),
			out2               => s_out2(1,16),
			lock_lower_row_out => s_locks_lower_out(1,16),
			lock_lower_row_in  => s_locks_lower_in(1,16),
			in1                => s_in1(1,16),
			in2                => s_in2(1,16),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(16)
		);
	s_in1(1,16)            <= s_out1(2,16);
	s_in2(1,16)            <= s_out2(2,17);
	s_locks_lower_in(1,16) <= s_locks_lower_out(2,16);

		normal_cell_1_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,17),
			fetch              => s_fetch(1,17),
			data_in            => s_data_in(1,17),
			data_out           => s_data_out(1,17),
			out1               => s_out1(1,17),
			out2               => s_out2(1,17),
			lock_lower_row_out => s_locks_lower_out(1,17),
			lock_lower_row_in  => s_locks_lower_in(1,17),
			in1                => s_in1(1,17),
			in2                => s_in2(1,17),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(17)
		);
	s_in1(1,17)            <= s_out1(2,17);
	s_in2(1,17)            <= s_out2(2,18);
	s_locks_lower_in(1,17) <= s_locks_lower_out(2,17);

		normal_cell_1_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,18),
			fetch              => s_fetch(1,18),
			data_in            => s_data_in(1,18),
			data_out           => s_data_out(1,18),
			out1               => s_out1(1,18),
			out2               => s_out2(1,18),
			lock_lower_row_out => s_locks_lower_out(1,18),
			lock_lower_row_in  => s_locks_lower_in(1,18),
			in1                => s_in1(1,18),
			in2                => s_in2(1,18),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(18)
		);
	s_in1(1,18)            <= s_out1(2,18);
	s_in2(1,18)            <= s_out2(2,19);
	s_locks_lower_in(1,18) <= s_locks_lower_out(2,18);

		normal_cell_1_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,19),
			fetch              => s_fetch(1,19),
			data_in            => s_data_in(1,19),
			data_out           => s_data_out(1,19),
			out1               => s_out1(1,19),
			out2               => s_out2(1,19),
			lock_lower_row_out => s_locks_lower_out(1,19),
			lock_lower_row_in  => s_locks_lower_in(1,19),
			in1                => s_in1(1,19),
			in2                => s_in2(1,19),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(19)
		);
	s_in1(1,19)            <= s_out1(2,19);
	s_in2(1,19)            <= s_out2(2,20);
	s_locks_lower_in(1,19) <= s_locks_lower_out(2,19);

		normal_cell_1_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,20),
			fetch              => s_fetch(1,20),
			data_in            => s_data_in(1,20),
			data_out           => s_data_out(1,20),
			out1               => s_out1(1,20),
			out2               => s_out2(1,20),
			lock_lower_row_out => s_locks_lower_out(1,20),
			lock_lower_row_in  => s_locks_lower_in(1,20),
			in1                => s_in1(1,20),
			in2                => s_in2(1,20),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(20)
		);
	s_in1(1,20)            <= s_out1(2,20);
	s_in2(1,20)            <= s_out2(2,21);
	s_locks_lower_in(1,20) <= s_locks_lower_out(2,20);

		normal_cell_1_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,21),
			fetch              => s_fetch(1,21),
			data_in            => s_data_in(1,21),
			data_out           => s_data_out(1,21),
			out1               => s_out1(1,21),
			out2               => s_out2(1,21),
			lock_lower_row_out => s_locks_lower_out(1,21),
			lock_lower_row_in  => s_locks_lower_in(1,21),
			in1                => s_in1(1,21),
			in2                => s_in2(1,21),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(21)
		);
	s_in1(1,21)            <= s_out1(2,21);
	s_in2(1,21)            <= s_out2(2,22);
	s_locks_lower_in(1,21) <= s_locks_lower_out(2,21);

		normal_cell_1_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,22),
			fetch              => s_fetch(1,22),
			data_in            => s_data_in(1,22),
			data_out           => s_data_out(1,22),
			out1               => s_out1(1,22),
			out2               => s_out2(1,22),
			lock_lower_row_out => s_locks_lower_out(1,22),
			lock_lower_row_in  => s_locks_lower_in(1,22),
			in1                => s_in1(1,22),
			in2                => s_in2(1,22),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(22)
		);
	s_in1(1,22)            <= s_out1(2,22);
	s_in2(1,22)            <= s_out2(2,23);
	s_locks_lower_in(1,22) <= s_locks_lower_out(2,22);

		normal_cell_1_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,23),
			fetch              => s_fetch(1,23),
			data_in            => s_data_in(1,23),
			data_out           => s_data_out(1,23),
			out1               => s_out1(1,23),
			out2               => s_out2(1,23),
			lock_lower_row_out => s_locks_lower_out(1,23),
			lock_lower_row_in  => s_locks_lower_in(1,23),
			in1                => s_in1(1,23),
			in2                => s_in2(1,23),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(23)
		);
	s_in1(1,23)            <= s_out1(2,23);
	s_in2(1,23)            <= s_out2(2,24);
	s_locks_lower_in(1,23) <= s_locks_lower_out(2,23);

		normal_cell_1_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,24),
			fetch              => s_fetch(1,24),
			data_in            => s_data_in(1,24),
			data_out           => s_data_out(1,24),
			out1               => s_out1(1,24),
			out2               => s_out2(1,24),
			lock_lower_row_out => s_locks_lower_out(1,24),
			lock_lower_row_in  => s_locks_lower_in(1,24),
			in1                => s_in1(1,24),
			in2                => s_in2(1,24),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(24)
		);
	s_in1(1,24)            <= s_out1(2,24);
	s_in2(1,24)            <= s_out2(2,25);
	s_locks_lower_in(1,24) <= s_locks_lower_out(2,24);

		normal_cell_1_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,25),
			fetch              => s_fetch(1,25),
			data_in            => s_data_in(1,25),
			data_out           => s_data_out(1,25),
			out1               => s_out1(1,25),
			out2               => s_out2(1,25),
			lock_lower_row_out => s_locks_lower_out(1,25),
			lock_lower_row_in  => s_locks_lower_in(1,25),
			in1                => s_in1(1,25),
			in2                => s_in2(1,25),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(25)
		);
	s_in1(1,25)            <= s_out1(2,25);
	s_in2(1,25)            <= s_out2(2,26);
	s_locks_lower_in(1,25) <= s_locks_lower_out(2,25);

		normal_cell_1_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,26),
			fetch              => s_fetch(1,26),
			data_in            => s_data_in(1,26),
			data_out           => s_data_out(1,26),
			out1               => s_out1(1,26),
			out2               => s_out2(1,26),
			lock_lower_row_out => s_locks_lower_out(1,26),
			lock_lower_row_in  => s_locks_lower_in(1,26),
			in1                => s_in1(1,26),
			in2                => s_in2(1,26),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(26)
		);
	s_in1(1,26)            <= s_out1(2,26);
	s_in2(1,26)            <= s_out2(2,27);
	s_locks_lower_in(1,26) <= s_locks_lower_out(2,26);

		normal_cell_1_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,27),
			fetch              => s_fetch(1,27),
			data_in            => s_data_in(1,27),
			data_out           => s_data_out(1,27),
			out1               => s_out1(1,27),
			out2               => s_out2(1,27),
			lock_lower_row_out => s_locks_lower_out(1,27),
			lock_lower_row_in  => s_locks_lower_in(1,27),
			in1                => s_in1(1,27),
			in2                => s_in2(1,27),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(27)
		);
	s_in1(1,27)            <= s_out1(2,27);
	s_in2(1,27)            <= s_out2(2,28);
	s_locks_lower_in(1,27) <= s_locks_lower_out(2,27);

		normal_cell_1_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,28),
			fetch              => s_fetch(1,28),
			data_in            => s_data_in(1,28),
			data_out           => s_data_out(1,28),
			out1               => s_out1(1,28),
			out2               => s_out2(1,28),
			lock_lower_row_out => s_locks_lower_out(1,28),
			lock_lower_row_in  => s_locks_lower_in(1,28),
			in1                => s_in1(1,28),
			in2                => s_in2(1,28),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(28)
		);
	s_in1(1,28)            <= s_out1(2,28);
	s_in2(1,28)            <= s_out2(2,29);
	s_locks_lower_in(1,28) <= s_locks_lower_out(2,28);

		normal_cell_1_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,29),
			fetch              => s_fetch(1,29),
			data_in            => s_data_in(1,29),
			data_out           => s_data_out(1,29),
			out1               => s_out1(1,29),
			out2               => s_out2(1,29),
			lock_lower_row_out => s_locks_lower_out(1,29),
			lock_lower_row_in  => s_locks_lower_in(1,29),
			in1                => s_in1(1,29),
			in2                => s_in2(1,29),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(29)
		);
	s_in1(1,29)            <= s_out1(2,29);
	s_in2(1,29)            <= s_out2(2,30);
	s_locks_lower_in(1,29) <= s_locks_lower_out(2,29);

		normal_cell_1_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,30),
			fetch              => s_fetch(1,30),
			data_in            => s_data_in(1,30),
			data_out           => s_data_out(1,30),
			out1               => s_out1(1,30),
			out2               => s_out2(1,30),
			lock_lower_row_out => s_locks_lower_out(1,30),
			lock_lower_row_in  => s_locks_lower_in(1,30),
			in1                => s_in1(1,30),
			in2                => s_in2(1,30),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(30)
		);
	s_in1(1,30)            <= s_out1(2,30);
	s_in2(1,30)            <= s_out2(2,31);
	s_locks_lower_in(1,30) <= s_locks_lower_out(2,30);

		normal_cell_1_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,31),
			fetch              => s_fetch(1,31),
			data_in            => s_data_in(1,31),
			data_out           => s_data_out(1,31),
			out1               => s_out1(1,31),
			out2               => s_out2(1,31),
			lock_lower_row_out => s_locks_lower_out(1,31),
			lock_lower_row_in  => s_locks_lower_in(1,31),
			in1                => s_in1(1,31),
			in2                => s_in2(1,31),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(31)
		);
	s_in1(1,31)            <= s_out1(2,31);
	s_in2(1,31)            <= s_out2(2,32);
	s_locks_lower_in(1,31) <= s_locks_lower_out(2,31);

		normal_cell_1_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,32),
			fetch              => s_fetch(1,32),
			data_in            => s_data_in(1,32),
			data_out           => s_data_out(1,32),
			out1               => s_out1(1,32),
			out2               => s_out2(1,32),
			lock_lower_row_out => s_locks_lower_out(1,32),
			lock_lower_row_in  => s_locks_lower_in(1,32),
			in1                => s_in1(1,32),
			in2                => s_in2(1,32),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(32)
		);
	s_in1(1,32)            <= s_out1(2,32);
	s_in2(1,32)            <= s_out2(2,33);
	s_locks_lower_in(1,32) <= s_locks_lower_out(2,32);

		normal_cell_1_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,33),
			fetch              => s_fetch(1,33),
			data_in            => s_data_in(1,33),
			data_out           => s_data_out(1,33),
			out1               => s_out1(1,33),
			out2               => s_out2(1,33),
			lock_lower_row_out => s_locks_lower_out(1,33),
			lock_lower_row_in  => s_locks_lower_in(1,33),
			in1                => s_in1(1,33),
			in2                => s_in2(1,33),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(33)
		);
	s_in1(1,33)            <= s_out1(2,33);
	s_in2(1,33)            <= s_out2(2,34);
	s_locks_lower_in(1,33) <= s_locks_lower_out(2,33);

		normal_cell_1_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,34),
			fetch              => s_fetch(1,34),
			data_in            => s_data_in(1,34),
			data_out           => s_data_out(1,34),
			out1               => s_out1(1,34),
			out2               => s_out2(1,34),
			lock_lower_row_out => s_locks_lower_out(1,34),
			lock_lower_row_in  => s_locks_lower_in(1,34),
			in1                => s_in1(1,34),
			in2                => s_in2(1,34),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(34)
		);
	s_in1(1,34)            <= s_out1(2,34);
	s_in2(1,34)            <= s_out2(2,35);
	s_locks_lower_in(1,34) <= s_locks_lower_out(2,34);

		normal_cell_1_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,35),
			fetch              => s_fetch(1,35),
			data_in            => s_data_in(1,35),
			data_out           => s_data_out(1,35),
			out1               => s_out1(1,35),
			out2               => s_out2(1,35),
			lock_lower_row_out => s_locks_lower_out(1,35),
			lock_lower_row_in  => s_locks_lower_in(1,35),
			in1                => s_in1(1,35),
			in2                => s_in2(1,35),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(35)
		);
	s_in1(1,35)            <= s_out1(2,35);
	s_in2(1,35)            <= s_out2(2,36);
	s_locks_lower_in(1,35) <= s_locks_lower_out(2,35);

		normal_cell_1_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,36),
			fetch              => s_fetch(1,36),
			data_in            => s_data_in(1,36),
			data_out           => s_data_out(1,36),
			out1               => s_out1(1,36),
			out2               => s_out2(1,36),
			lock_lower_row_out => s_locks_lower_out(1,36),
			lock_lower_row_in  => s_locks_lower_in(1,36),
			in1                => s_in1(1,36),
			in2                => s_in2(1,36),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(36)
		);
	s_in1(1,36)            <= s_out1(2,36);
	s_in2(1,36)            <= s_out2(2,37);
	s_locks_lower_in(1,36) <= s_locks_lower_out(2,36);

		normal_cell_1_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,37),
			fetch              => s_fetch(1,37),
			data_in            => s_data_in(1,37),
			data_out           => s_data_out(1,37),
			out1               => s_out1(1,37),
			out2               => s_out2(1,37),
			lock_lower_row_out => s_locks_lower_out(1,37),
			lock_lower_row_in  => s_locks_lower_in(1,37),
			in1                => s_in1(1,37),
			in2                => s_in2(1,37),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(37)
		);
	s_in1(1,37)            <= s_out1(2,37);
	s_in2(1,37)            <= s_out2(2,38);
	s_locks_lower_in(1,37) <= s_locks_lower_out(2,37);

		normal_cell_1_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,38),
			fetch              => s_fetch(1,38),
			data_in            => s_data_in(1,38),
			data_out           => s_data_out(1,38),
			out1               => s_out1(1,38),
			out2               => s_out2(1,38),
			lock_lower_row_out => s_locks_lower_out(1,38),
			lock_lower_row_in  => s_locks_lower_in(1,38),
			in1                => s_in1(1,38),
			in2                => s_in2(1,38),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(38)
		);
	s_in1(1,38)            <= s_out1(2,38);
	s_in2(1,38)            <= s_out2(2,39);
	s_locks_lower_in(1,38) <= s_locks_lower_out(2,38);

		normal_cell_1_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,39),
			fetch              => s_fetch(1,39),
			data_in            => s_data_in(1,39),
			data_out           => s_data_out(1,39),
			out1               => s_out1(1,39),
			out2               => s_out2(1,39),
			lock_lower_row_out => s_locks_lower_out(1,39),
			lock_lower_row_in  => s_locks_lower_in(1,39),
			in1                => s_in1(1,39),
			in2                => s_in2(1,39),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(39)
		);
	s_in1(1,39)            <= s_out1(2,39);
	s_in2(1,39)            <= s_out2(2,40);
	s_locks_lower_in(1,39) <= s_locks_lower_out(2,39);

		normal_cell_1_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,40),
			fetch              => s_fetch(1,40),
			data_in            => s_data_in(1,40),
			data_out           => s_data_out(1,40),
			out1               => s_out1(1,40),
			out2               => s_out2(1,40),
			lock_lower_row_out => s_locks_lower_out(1,40),
			lock_lower_row_in  => s_locks_lower_in(1,40),
			in1                => s_in1(1,40),
			in2                => s_in2(1,40),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(40)
		);
	s_in1(1,40)            <= s_out1(2,40);
	s_in2(1,40)            <= s_out2(2,41);
	s_locks_lower_in(1,40) <= s_locks_lower_out(2,40);

		normal_cell_1_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,41),
			fetch              => s_fetch(1,41),
			data_in            => s_data_in(1,41),
			data_out           => s_data_out(1,41),
			out1               => s_out1(1,41),
			out2               => s_out2(1,41),
			lock_lower_row_out => s_locks_lower_out(1,41),
			lock_lower_row_in  => s_locks_lower_in(1,41),
			in1                => s_in1(1,41),
			in2                => s_in2(1,41),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(41)
		);
	s_in1(1,41)            <= s_out1(2,41);
	s_in2(1,41)            <= s_out2(2,42);
	s_locks_lower_in(1,41) <= s_locks_lower_out(2,41);

		normal_cell_1_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,42),
			fetch              => s_fetch(1,42),
			data_in            => s_data_in(1,42),
			data_out           => s_data_out(1,42),
			out1               => s_out1(1,42),
			out2               => s_out2(1,42),
			lock_lower_row_out => s_locks_lower_out(1,42),
			lock_lower_row_in  => s_locks_lower_in(1,42),
			in1                => s_in1(1,42),
			in2                => s_in2(1,42),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(42)
		);
	s_in1(1,42)            <= s_out1(2,42);
	s_in2(1,42)            <= s_out2(2,43);
	s_locks_lower_in(1,42) <= s_locks_lower_out(2,42);

		normal_cell_1_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,43),
			fetch              => s_fetch(1,43),
			data_in            => s_data_in(1,43),
			data_out           => s_data_out(1,43),
			out1               => s_out1(1,43),
			out2               => s_out2(1,43),
			lock_lower_row_out => s_locks_lower_out(1,43),
			lock_lower_row_in  => s_locks_lower_in(1,43),
			in1                => s_in1(1,43),
			in2                => s_in2(1,43),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(43)
		);
	s_in1(1,43)            <= s_out1(2,43);
	s_in2(1,43)            <= s_out2(2,44);
	s_locks_lower_in(1,43) <= s_locks_lower_out(2,43);

		normal_cell_1_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,44),
			fetch              => s_fetch(1,44),
			data_in            => s_data_in(1,44),
			data_out           => s_data_out(1,44),
			out1               => s_out1(1,44),
			out2               => s_out2(1,44),
			lock_lower_row_out => s_locks_lower_out(1,44),
			lock_lower_row_in  => s_locks_lower_in(1,44),
			in1                => s_in1(1,44),
			in2                => s_in2(1,44),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(44)
		);
	s_in1(1,44)            <= s_out1(2,44);
	s_in2(1,44)            <= s_out2(2,45);
	s_locks_lower_in(1,44) <= s_locks_lower_out(2,44);

		normal_cell_1_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,45),
			fetch              => s_fetch(1,45),
			data_in            => s_data_in(1,45),
			data_out           => s_data_out(1,45),
			out1               => s_out1(1,45),
			out2               => s_out2(1,45),
			lock_lower_row_out => s_locks_lower_out(1,45),
			lock_lower_row_in  => s_locks_lower_in(1,45),
			in1                => s_in1(1,45),
			in2                => s_in2(1,45),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(45)
		);
	s_in1(1,45)            <= s_out1(2,45);
	s_in2(1,45)            <= s_out2(2,46);
	s_locks_lower_in(1,45) <= s_locks_lower_out(2,45);

		normal_cell_1_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,46),
			fetch              => s_fetch(1,46),
			data_in            => s_data_in(1,46),
			data_out           => s_data_out(1,46),
			out1               => s_out1(1,46),
			out2               => s_out2(1,46),
			lock_lower_row_out => s_locks_lower_out(1,46),
			lock_lower_row_in  => s_locks_lower_in(1,46),
			in1                => s_in1(1,46),
			in2                => s_in2(1,46),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(46)
		);
	s_in1(1,46)            <= s_out1(2,46);
	s_in2(1,46)            <= s_out2(2,47);
	s_locks_lower_in(1,46) <= s_locks_lower_out(2,46);

		normal_cell_1_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,47),
			fetch              => s_fetch(1,47),
			data_in            => s_data_in(1,47),
			data_out           => s_data_out(1,47),
			out1               => s_out1(1,47),
			out2               => s_out2(1,47),
			lock_lower_row_out => s_locks_lower_out(1,47),
			lock_lower_row_in  => s_locks_lower_in(1,47),
			in1                => s_in1(1,47),
			in2                => s_in2(1,47),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(47)
		);
	s_in1(1,47)            <= s_out1(2,47);
	s_in2(1,47)            <= s_out2(2,48);
	s_locks_lower_in(1,47) <= s_locks_lower_out(2,47);

		normal_cell_1_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,48),
			fetch              => s_fetch(1,48),
			data_in            => s_data_in(1,48),
			data_out           => s_data_out(1,48),
			out1               => s_out1(1,48),
			out2               => s_out2(1,48),
			lock_lower_row_out => s_locks_lower_out(1,48),
			lock_lower_row_in  => s_locks_lower_in(1,48),
			in1                => s_in1(1,48),
			in2                => s_in2(1,48),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(48)
		);
	s_in1(1,48)            <= s_out1(2,48);
	s_in2(1,48)            <= s_out2(2,49);
	s_locks_lower_in(1,48) <= s_locks_lower_out(2,48);

		normal_cell_1_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,49),
			fetch              => s_fetch(1,49),
			data_in            => s_data_in(1,49),
			data_out           => s_data_out(1,49),
			out1               => s_out1(1,49),
			out2               => s_out2(1,49),
			lock_lower_row_out => s_locks_lower_out(1,49),
			lock_lower_row_in  => s_locks_lower_in(1,49),
			in1                => s_in1(1,49),
			in2                => s_in2(1,49),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(49)
		);
	s_in1(1,49)            <= s_out1(2,49);
	s_in2(1,49)            <= s_out2(2,50);
	s_locks_lower_in(1,49) <= s_locks_lower_out(2,49);

		normal_cell_1_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,50),
			fetch              => s_fetch(1,50),
			data_in            => s_data_in(1,50),
			data_out           => s_data_out(1,50),
			out1               => s_out1(1,50),
			out2               => s_out2(1,50),
			lock_lower_row_out => s_locks_lower_out(1,50),
			lock_lower_row_in  => s_locks_lower_in(1,50),
			in1                => s_in1(1,50),
			in2                => s_in2(1,50),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(50)
		);
	s_in1(1,50)            <= s_out1(2,50);
	s_in2(1,50)            <= s_out2(2,51);
	s_locks_lower_in(1,50) <= s_locks_lower_out(2,50);

		normal_cell_1_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,51),
			fetch              => s_fetch(1,51),
			data_in            => s_data_in(1,51),
			data_out           => s_data_out(1,51),
			out1               => s_out1(1,51),
			out2               => s_out2(1,51),
			lock_lower_row_out => s_locks_lower_out(1,51),
			lock_lower_row_in  => s_locks_lower_in(1,51),
			in1                => s_in1(1,51),
			in2                => s_in2(1,51),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(51)
		);
	s_in1(1,51)            <= s_out1(2,51);
	s_in2(1,51)            <= s_out2(2,52);
	s_locks_lower_in(1,51) <= s_locks_lower_out(2,51);

		normal_cell_1_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,52),
			fetch              => s_fetch(1,52),
			data_in            => s_data_in(1,52),
			data_out           => s_data_out(1,52),
			out1               => s_out1(1,52),
			out2               => s_out2(1,52),
			lock_lower_row_out => s_locks_lower_out(1,52),
			lock_lower_row_in  => s_locks_lower_in(1,52),
			in1                => s_in1(1,52),
			in2                => s_in2(1,52),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(52)
		);
	s_in1(1,52)            <= s_out1(2,52);
	s_in2(1,52)            <= s_out2(2,53);
	s_locks_lower_in(1,52) <= s_locks_lower_out(2,52);

		normal_cell_1_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,53),
			fetch              => s_fetch(1,53),
			data_in            => s_data_in(1,53),
			data_out           => s_data_out(1,53),
			out1               => s_out1(1,53),
			out2               => s_out2(1,53),
			lock_lower_row_out => s_locks_lower_out(1,53),
			lock_lower_row_in  => s_locks_lower_in(1,53),
			in1                => s_in1(1,53),
			in2                => s_in2(1,53),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(53)
		);
	s_in1(1,53)            <= s_out1(2,53);
	s_in2(1,53)            <= s_out2(2,54);
	s_locks_lower_in(1,53) <= s_locks_lower_out(2,53);

		normal_cell_1_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,54),
			fetch              => s_fetch(1,54),
			data_in            => s_data_in(1,54),
			data_out           => s_data_out(1,54),
			out1               => s_out1(1,54),
			out2               => s_out2(1,54),
			lock_lower_row_out => s_locks_lower_out(1,54),
			lock_lower_row_in  => s_locks_lower_in(1,54),
			in1                => s_in1(1,54),
			in2                => s_in2(1,54),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(54)
		);
	s_in1(1,54)            <= s_out1(2,54);
	s_in2(1,54)            <= s_out2(2,55);
	s_locks_lower_in(1,54) <= s_locks_lower_out(2,54);

		normal_cell_1_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,55),
			fetch              => s_fetch(1,55),
			data_in            => s_data_in(1,55),
			data_out           => s_data_out(1,55),
			out1               => s_out1(1,55),
			out2               => s_out2(1,55),
			lock_lower_row_out => s_locks_lower_out(1,55),
			lock_lower_row_in  => s_locks_lower_in(1,55),
			in1                => s_in1(1,55),
			in2                => s_in2(1,55),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(55)
		);
	s_in1(1,55)            <= s_out1(2,55);
	s_in2(1,55)            <= s_out2(2,56);
	s_locks_lower_in(1,55) <= s_locks_lower_out(2,55);

		normal_cell_1_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,56),
			fetch              => s_fetch(1,56),
			data_in            => s_data_in(1,56),
			data_out           => s_data_out(1,56),
			out1               => s_out1(1,56),
			out2               => s_out2(1,56),
			lock_lower_row_out => s_locks_lower_out(1,56),
			lock_lower_row_in  => s_locks_lower_in(1,56),
			in1                => s_in1(1,56),
			in2                => s_in2(1,56),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(56)
		);
	s_in1(1,56)            <= s_out1(2,56);
	s_in2(1,56)            <= s_out2(2,57);
	s_locks_lower_in(1,56) <= s_locks_lower_out(2,56);

		normal_cell_1_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,57),
			fetch              => s_fetch(1,57),
			data_in            => s_data_in(1,57),
			data_out           => s_data_out(1,57),
			out1               => s_out1(1,57),
			out2               => s_out2(1,57),
			lock_lower_row_out => s_locks_lower_out(1,57),
			lock_lower_row_in  => s_locks_lower_in(1,57),
			in1                => s_in1(1,57),
			in2                => s_in2(1,57),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(57)
		);
	s_in1(1,57)            <= s_out1(2,57);
	s_in2(1,57)            <= s_out2(2,58);
	s_locks_lower_in(1,57) <= s_locks_lower_out(2,57);

		normal_cell_1_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,58),
			fetch              => s_fetch(1,58),
			data_in            => s_data_in(1,58),
			data_out           => s_data_out(1,58),
			out1               => s_out1(1,58),
			out2               => s_out2(1,58),
			lock_lower_row_out => s_locks_lower_out(1,58),
			lock_lower_row_in  => s_locks_lower_in(1,58),
			in1                => s_in1(1,58),
			in2                => s_in2(1,58),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(58)
		);
	s_in1(1,58)            <= s_out1(2,58);
	s_in2(1,58)            <= s_out2(2,59);
	s_locks_lower_in(1,58) <= s_locks_lower_out(2,58);

		normal_cell_1_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,59),
			fetch              => s_fetch(1,59),
			data_in            => s_data_in(1,59),
			data_out           => s_data_out(1,59),
			out1               => s_out1(1,59),
			out2               => s_out2(1,59),
			lock_lower_row_out => s_locks_lower_out(1,59),
			lock_lower_row_in  => s_locks_lower_in(1,59),
			in1                => s_in1(1,59),
			in2                => s_in2(1,59),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(59)
		);
	s_in1(1,59)            <= s_out1(2,59);
	s_in2(1,59)            <= s_out2(2,60);
	s_locks_lower_in(1,59) <= s_locks_lower_out(2,59);

		last_col_cell_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(1,60),
			fetch              => s_fetch(1,60),
			data_in            => s_data_in(1,60),
			data_out           => s_data_out(1,60),
			out1               => s_out1(1,60),
			out2               => s_out2(1,60),
			lock_lower_row_out => s_locks_lower_out(1,60),
			lock_lower_row_in  => s_locks_lower_in(1,60),
			in1                => s_in1(1,60),
			in2                => (others => '0'),
			lock_row           => s_locks(1),
			piv_found          => s_piv_found,
			row_data           => s_row_data(1),
			col_data           => s_col_data(60)
		);
	s_in1(1,60)            <= s_out1(2,60);
	s_locks_lower_in(1,60) <= s_locks_lower_out(2,60);

		normal_cell_2_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,1),
			fetch              => s_fetch(2,1),
			data_in            => s_data_in(2,1),
			data_out           => s_data_out(2,1),
			out1               => s_out1(2,1),
			out2               => s_out2(2,1),
			lock_lower_row_out => s_locks_lower_out(2,1),
			lock_lower_row_in  => s_locks_lower_in(2,1),
			in1                => s_in1(2,1),
			in2                => s_in2(2,1),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(1)
		);
	s_in1(2,1)            <= s_out1(3,1);
	s_in2(2,1)            <= s_out2(3,2);
	s_locks_lower_in(2,1) <= s_locks_lower_out(3,1);

		normal_cell_2_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,2),
			fetch              => s_fetch(2,2),
			data_in            => s_data_in(2,2),
			data_out           => s_data_out(2,2),
			out1               => s_out1(2,2),
			out2               => s_out2(2,2),
			lock_lower_row_out => s_locks_lower_out(2,2),
			lock_lower_row_in  => s_locks_lower_in(2,2),
			in1                => s_in1(2,2),
			in2                => s_in2(2,2),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(2)
		);
	s_in1(2,2)            <= s_out1(3,2);
	s_in2(2,2)            <= s_out2(3,3);
	s_locks_lower_in(2,2) <= s_locks_lower_out(3,2);

		normal_cell_2_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,3),
			fetch              => s_fetch(2,3),
			data_in            => s_data_in(2,3),
			data_out           => s_data_out(2,3),
			out1               => s_out1(2,3),
			out2               => s_out2(2,3),
			lock_lower_row_out => s_locks_lower_out(2,3),
			lock_lower_row_in  => s_locks_lower_in(2,3),
			in1                => s_in1(2,3),
			in2                => s_in2(2,3),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(3)
		);
	s_in1(2,3)            <= s_out1(3,3);
	s_in2(2,3)            <= s_out2(3,4);
	s_locks_lower_in(2,3) <= s_locks_lower_out(3,3);

		normal_cell_2_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,4),
			fetch              => s_fetch(2,4),
			data_in            => s_data_in(2,4),
			data_out           => s_data_out(2,4),
			out1               => s_out1(2,4),
			out2               => s_out2(2,4),
			lock_lower_row_out => s_locks_lower_out(2,4),
			lock_lower_row_in  => s_locks_lower_in(2,4),
			in1                => s_in1(2,4),
			in2                => s_in2(2,4),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(4)
		);
	s_in1(2,4)            <= s_out1(3,4);
	s_in2(2,4)            <= s_out2(3,5);
	s_locks_lower_in(2,4) <= s_locks_lower_out(3,4);

		normal_cell_2_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,5),
			fetch              => s_fetch(2,5),
			data_in            => s_data_in(2,5),
			data_out           => s_data_out(2,5),
			out1               => s_out1(2,5),
			out2               => s_out2(2,5),
			lock_lower_row_out => s_locks_lower_out(2,5),
			lock_lower_row_in  => s_locks_lower_in(2,5),
			in1                => s_in1(2,5),
			in2                => s_in2(2,5),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(5)
		);
	s_in1(2,5)            <= s_out1(3,5);
	s_in2(2,5)            <= s_out2(3,6);
	s_locks_lower_in(2,5) <= s_locks_lower_out(3,5);

		normal_cell_2_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,6),
			fetch              => s_fetch(2,6),
			data_in            => s_data_in(2,6),
			data_out           => s_data_out(2,6),
			out1               => s_out1(2,6),
			out2               => s_out2(2,6),
			lock_lower_row_out => s_locks_lower_out(2,6),
			lock_lower_row_in  => s_locks_lower_in(2,6),
			in1                => s_in1(2,6),
			in2                => s_in2(2,6),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(6)
		);
	s_in1(2,6)            <= s_out1(3,6);
	s_in2(2,6)            <= s_out2(3,7);
	s_locks_lower_in(2,6) <= s_locks_lower_out(3,6);

		normal_cell_2_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,7),
			fetch              => s_fetch(2,7),
			data_in            => s_data_in(2,7),
			data_out           => s_data_out(2,7),
			out1               => s_out1(2,7),
			out2               => s_out2(2,7),
			lock_lower_row_out => s_locks_lower_out(2,7),
			lock_lower_row_in  => s_locks_lower_in(2,7),
			in1                => s_in1(2,7),
			in2                => s_in2(2,7),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(7)
		);
	s_in1(2,7)            <= s_out1(3,7);
	s_in2(2,7)            <= s_out2(3,8);
	s_locks_lower_in(2,7) <= s_locks_lower_out(3,7);

		normal_cell_2_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,8),
			fetch              => s_fetch(2,8),
			data_in            => s_data_in(2,8),
			data_out           => s_data_out(2,8),
			out1               => s_out1(2,8),
			out2               => s_out2(2,8),
			lock_lower_row_out => s_locks_lower_out(2,8),
			lock_lower_row_in  => s_locks_lower_in(2,8),
			in1                => s_in1(2,8),
			in2                => s_in2(2,8),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(8)
		);
	s_in1(2,8)            <= s_out1(3,8);
	s_in2(2,8)            <= s_out2(3,9);
	s_locks_lower_in(2,8) <= s_locks_lower_out(3,8);

		normal_cell_2_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,9),
			fetch              => s_fetch(2,9),
			data_in            => s_data_in(2,9),
			data_out           => s_data_out(2,9),
			out1               => s_out1(2,9),
			out2               => s_out2(2,9),
			lock_lower_row_out => s_locks_lower_out(2,9),
			lock_lower_row_in  => s_locks_lower_in(2,9),
			in1                => s_in1(2,9),
			in2                => s_in2(2,9),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(9)
		);
	s_in1(2,9)            <= s_out1(3,9);
	s_in2(2,9)            <= s_out2(3,10);
	s_locks_lower_in(2,9) <= s_locks_lower_out(3,9);

		normal_cell_2_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,10),
			fetch              => s_fetch(2,10),
			data_in            => s_data_in(2,10),
			data_out           => s_data_out(2,10),
			out1               => s_out1(2,10),
			out2               => s_out2(2,10),
			lock_lower_row_out => s_locks_lower_out(2,10),
			lock_lower_row_in  => s_locks_lower_in(2,10),
			in1                => s_in1(2,10),
			in2                => s_in2(2,10),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(10)
		);
	s_in1(2,10)            <= s_out1(3,10);
	s_in2(2,10)            <= s_out2(3,11);
	s_locks_lower_in(2,10) <= s_locks_lower_out(3,10);

		normal_cell_2_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,11),
			fetch              => s_fetch(2,11),
			data_in            => s_data_in(2,11),
			data_out           => s_data_out(2,11),
			out1               => s_out1(2,11),
			out2               => s_out2(2,11),
			lock_lower_row_out => s_locks_lower_out(2,11),
			lock_lower_row_in  => s_locks_lower_in(2,11),
			in1                => s_in1(2,11),
			in2                => s_in2(2,11),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(11)
		);
	s_in1(2,11)            <= s_out1(3,11);
	s_in2(2,11)            <= s_out2(3,12);
	s_locks_lower_in(2,11) <= s_locks_lower_out(3,11);

		normal_cell_2_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,12),
			fetch              => s_fetch(2,12),
			data_in            => s_data_in(2,12),
			data_out           => s_data_out(2,12),
			out1               => s_out1(2,12),
			out2               => s_out2(2,12),
			lock_lower_row_out => s_locks_lower_out(2,12),
			lock_lower_row_in  => s_locks_lower_in(2,12),
			in1                => s_in1(2,12),
			in2                => s_in2(2,12),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(12)
		);
	s_in1(2,12)            <= s_out1(3,12);
	s_in2(2,12)            <= s_out2(3,13);
	s_locks_lower_in(2,12) <= s_locks_lower_out(3,12);

		normal_cell_2_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,13),
			fetch              => s_fetch(2,13),
			data_in            => s_data_in(2,13),
			data_out           => s_data_out(2,13),
			out1               => s_out1(2,13),
			out2               => s_out2(2,13),
			lock_lower_row_out => s_locks_lower_out(2,13),
			lock_lower_row_in  => s_locks_lower_in(2,13),
			in1                => s_in1(2,13),
			in2                => s_in2(2,13),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(13)
		);
	s_in1(2,13)            <= s_out1(3,13);
	s_in2(2,13)            <= s_out2(3,14);
	s_locks_lower_in(2,13) <= s_locks_lower_out(3,13);

		normal_cell_2_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,14),
			fetch              => s_fetch(2,14),
			data_in            => s_data_in(2,14),
			data_out           => s_data_out(2,14),
			out1               => s_out1(2,14),
			out2               => s_out2(2,14),
			lock_lower_row_out => s_locks_lower_out(2,14),
			lock_lower_row_in  => s_locks_lower_in(2,14),
			in1                => s_in1(2,14),
			in2                => s_in2(2,14),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(14)
		);
	s_in1(2,14)            <= s_out1(3,14);
	s_in2(2,14)            <= s_out2(3,15);
	s_locks_lower_in(2,14) <= s_locks_lower_out(3,14);

		normal_cell_2_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,15),
			fetch              => s_fetch(2,15),
			data_in            => s_data_in(2,15),
			data_out           => s_data_out(2,15),
			out1               => s_out1(2,15),
			out2               => s_out2(2,15),
			lock_lower_row_out => s_locks_lower_out(2,15),
			lock_lower_row_in  => s_locks_lower_in(2,15),
			in1                => s_in1(2,15),
			in2                => s_in2(2,15),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(15)
		);
	s_in1(2,15)            <= s_out1(3,15);
	s_in2(2,15)            <= s_out2(3,16);
	s_locks_lower_in(2,15) <= s_locks_lower_out(3,15);

		normal_cell_2_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,16),
			fetch              => s_fetch(2,16),
			data_in            => s_data_in(2,16),
			data_out           => s_data_out(2,16),
			out1               => s_out1(2,16),
			out2               => s_out2(2,16),
			lock_lower_row_out => s_locks_lower_out(2,16),
			lock_lower_row_in  => s_locks_lower_in(2,16),
			in1                => s_in1(2,16),
			in2                => s_in2(2,16),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(16)
		);
	s_in1(2,16)            <= s_out1(3,16);
	s_in2(2,16)            <= s_out2(3,17);
	s_locks_lower_in(2,16) <= s_locks_lower_out(3,16);

		normal_cell_2_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,17),
			fetch              => s_fetch(2,17),
			data_in            => s_data_in(2,17),
			data_out           => s_data_out(2,17),
			out1               => s_out1(2,17),
			out2               => s_out2(2,17),
			lock_lower_row_out => s_locks_lower_out(2,17),
			lock_lower_row_in  => s_locks_lower_in(2,17),
			in1                => s_in1(2,17),
			in2                => s_in2(2,17),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(17)
		);
	s_in1(2,17)            <= s_out1(3,17);
	s_in2(2,17)            <= s_out2(3,18);
	s_locks_lower_in(2,17) <= s_locks_lower_out(3,17);

		normal_cell_2_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,18),
			fetch              => s_fetch(2,18),
			data_in            => s_data_in(2,18),
			data_out           => s_data_out(2,18),
			out1               => s_out1(2,18),
			out2               => s_out2(2,18),
			lock_lower_row_out => s_locks_lower_out(2,18),
			lock_lower_row_in  => s_locks_lower_in(2,18),
			in1                => s_in1(2,18),
			in2                => s_in2(2,18),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(18)
		);
	s_in1(2,18)            <= s_out1(3,18);
	s_in2(2,18)            <= s_out2(3,19);
	s_locks_lower_in(2,18) <= s_locks_lower_out(3,18);

		normal_cell_2_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,19),
			fetch              => s_fetch(2,19),
			data_in            => s_data_in(2,19),
			data_out           => s_data_out(2,19),
			out1               => s_out1(2,19),
			out2               => s_out2(2,19),
			lock_lower_row_out => s_locks_lower_out(2,19),
			lock_lower_row_in  => s_locks_lower_in(2,19),
			in1                => s_in1(2,19),
			in2                => s_in2(2,19),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(19)
		);
	s_in1(2,19)            <= s_out1(3,19);
	s_in2(2,19)            <= s_out2(3,20);
	s_locks_lower_in(2,19) <= s_locks_lower_out(3,19);

		normal_cell_2_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,20),
			fetch              => s_fetch(2,20),
			data_in            => s_data_in(2,20),
			data_out           => s_data_out(2,20),
			out1               => s_out1(2,20),
			out2               => s_out2(2,20),
			lock_lower_row_out => s_locks_lower_out(2,20),
			lock_lower_row_in  => s_locks_lower_in(2,20),
			in1                => s_in1(2,20),
			in2                => s_in2(2,20),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(20)
		);
	s_in1(2,20)            <= s_out1(3,20);
	s_in2(2,20)            <= s_out2(3,21);
	s_locks_lower_in(2,20) <= s_locks_lower_out(3,20);

		normal_cell_2_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,21),
			fetch              => s_fetch(2,21),
			data_in            => s_data_in(2,21),
			data_out           => s_data_out(2,21),
			out1               => s_out1(2,21),
			out2               => s_out2(2,21),
			lock_lower_row_out => s_locks_lower_out(2,21),
			lock_lower_row_in  => s_locks_lower_in(2,21),
			in1                => s_in1(2,21),
			in2                => s_in2(2,21),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(21)
		);
	s_in1(2,21)            <= s_out1(3,21);
	s_in2(2,21)            <= s_out2(3,22);
	s_locks_lower_in(2,21) <= s_locks_lower_out(3,21);

		normal_cell_2_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,22),
			fetch              => s_fetch(2,22),
			data_in            => s_data_in(2,22),
			data_out           => s_data_out(2,22),
			out1               => s_out1(2,22),
			out2               => s_out2(2,22),
			lock_lower_row_out => s_locks_lower_out(2,22),
			lock_lower_row_in  => s_locks_lower_in(2,22),
			in1                => s_in1(2,22),
			in2                => s_in2(2,22),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(22)
		);
	s_in1(2,22)            <= s_out1(3,22);
	s_in2(2,22)            <= s_out2(3,23);
	s_locks_lower_in(2,22) <= s_locks_lower_out(3,22);

		normal_cell_2_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,23),
			fetch              => s_fetch(2,23),
			data_in            => s_data_in(2,23),
			data_out           => s_data_out(2,23),
			out1               => s_out1(2,23),
			out2               => s_out2(2,23),
			lock_lower_row_out => s_locks_lower_out(2,23),
			lock_lower_row_in  => s_locks_lower_in(2,23),
			in1                => s_in1(2,23),
			in2                => s_in2(2,23),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(23)
		);
	s_in1(2,23)            <= s_out1(3,23);
	s_in2(2,23)            <= s_out2(3,24);
	s_locks_lower_in(2,23) <= s_locks_lower_out(3,23);

		normal_cell_2_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,24),
			fetch              => s_fetch(2,24),
			data_in            => s_data_in(2,24),
			data_out           => s_data_out(2,24),
			out1               => s_out1(2,24),
			out2               => s_out2(2,24),
			lock_lower_row_out => s_locks_lower_out(2,24),
			lock_lower_row_in  => s_locks_lower_in(2,24),
			in1                => s_in1(2,24),
			in2                => s_in2(2,24),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(24)
		);
	s_in1(2,24)            <= s_out1(3,24);
	s_in2(2,24)            <= s_out2(3,25);
	s_locks_lower_in(2,24) <= s_locks_lower_out(3,24);

		normal_cell_2_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,25),
			fetch              => s_fetch(2,25),
			data_in            => s_data_in(2,25),
			data_out           => s_data_out(2,25),
			out1               => s_out1(2,25),
			out2               => s_out2(2,25),
			lock_lower_row_out => s_locks_lower_out(2,25),
			lock_lower_row_in  => s_locks_lower_in(2,25),
			in1                => s_in1(2,25),
			in2                => s_in2(2,25),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(25)
		);
	s_in1(2,25)            <= s_out1(3,25);
	s_in2(2,25)            <= s_out2(3,26);
	s_locks_lower_in(2,25) <= s_locks_lower_out(3,25);

		normal_cell_2_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,26),
			fetch              => s_fetch(2,26),
			data_in            => s_data_in(2,26),
			data_out           => s_data_out(2,26),
			out1               => s_out1(2,26),
			out2               => s_out2(2,26),
			lock_lower_row_out => s_locks_lower_out(2,26),
			lock_lower_row_in  => s_locks_lower_in(2,26),
			in1                => s_in1(2,26),
			in2                => s_in2(2,26),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(26)
		);
	s_in1(2,26)            <= s_out1(3,26);
	s_in2(2,26)            <= s_out2(3,27);
	s_locks_lower_in(2,26) <= s_locks_lower_out(3,26);

		normal_cell_2_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,27),
			fetch              => s_fetch(2,27),
			data_in            => s_data_in(2,27),
			data_out           => s_data_out(2,27),
			out1               => s_out1(2,27),
			out2               => s_out2(2,27),
			lock_lower_row_out => s_locks_lower_out(2,27),
			lock_lower_row_in  => s_locks_lower_in(2,27),
			in1                => s_in1(2,27),
			in2                => s_in2(2,27),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(27)
		);
	s_in1(2,27)            <= s_out1(3,27);
	s_in2(2,27)            <= s_out2(3,28);
	s_locks_lower_in(2,27) <= s_locks_lower_out(3,27);

		normal_cell_2_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,28),
			fetch              => s_fetch(2,28),
			data_in            => s_data_in(2,28),
			data_out           => s_data_out(2,28),
			out1               => s_out1(2,28),
			out2               => s_out2(2,28),
			lock_lower_row_out => s_locks_lower_out(2,28),
			lock_lower_row_in  => s_locks_lower_in(2,28),
			in1                => s_in1(2,28),
			in2                => s_in2(2,28),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(28)
		);
	s_in1(2,28)            <= s_out1(3,28);
	s_in2(2,28)            <= s_out2(3,29);
	s_locks_lower_in(2,28) <= s_locks_lower_out(3,28);

		normal_cell_2_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,29),
			fetch              => s_fetch(2,29),
			data_in            => s_data_in(2,29),
			data_out           => s_data_out(2,29),
			out1               => s_out1(2,29),
			out2               => s_out2(2,29),
			lock_lower_row_out => s_locks_lower_out(2,29),
			lock_lower_row_in  => s_locks_lower_in(2,29),
			in1                => s_in1(2,29),
			in2                => s_in2(2,29),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(29)
		);
	s_in1(2,29)            <= s_out1(3,29);
	s_in2(2,29)            <= s_out2(3,30);
	s_locks_lower_in(2,29) <= s_locks_lower_out(3,29);

		normal_cell_2_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,30),
			fetch              => s_fetch(2,30),
			data_in            => s_data_in(2,30),
			data_out           => s_data_out(2,30),
			out1               => s_out1(2,30),
			out2               => s_out2(2,30),
			lock_lower_row_out => s_locks_lower_out(2,30),
			lock_lower_row_in  => s_locks_lower_in(2,30),
			in1                => s_in1(2,30),
			in2                => s_in2(2,30),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(30)
		);
	s_in1(2,30)            <= s_out1(3,30);
	s_in2(2,30)            <= s_out2(3,31);
	s_locks_lower_in(2,30) <= s_locks_lower_out(3,30);

		normal_cell_2_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,31),
			fetch              => s_fetch(2,31),
			data_in            => s_data_in(2,31),
			data_out           => s_data_out(2,31),
			out1               => s_out1(2,31),
			out2               => s_out2(2,31),
			lock_lower_row_out => s_locks_lower_out(2,31),
			lock_lower_row_in  => s_locks_lower_in(2,31),
			in1                => s_in1(2,31),
			in2                => s_in2(2,31),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(31)
		);
	s_in1(2,31)            <= s_out1(3,31);
	s_in2(2,31)            <= s_out2(3,32);
	s_locks_lower_in(2,31) <= s_locks_lower_out(3,31);

		normal_cell_2_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,32),
			fetch              => s_fetch(2,32),
			data_in            => s_data_in(2,32),
			data_out           => s_data_out(2,32),
			out1               => s_out1(2,32),
			out2               => s_out2(2,32),
			lock_lower_row_out => s_locks_lower_out(2,32),
			lock_lower_row_in  => s_locks_lower_in(2,32),
			in1                => s_in1(2,32),
			in2                => s_in2(2,32),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(32)
		);
	s_in1(2,32)            <= s_out1(3,32);
	s_in2(2,32)            <= s_out2(3,33);
	s_locks_lower_in(2,32) <= s_locks_lower_out(3,32);

		normal_cell_2_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,33),
			fetch              => s_fetch(2,33),
			data_in            => s_data_in(2,33),
			data_out           => s_data_out(2,33),
			out1               => s_out1(2,33),
			out2               => s_out2(2,33),
			lock_lower_row_out => s_locks_lower_out(2,33),
			lock_lower_row_in  => s_locks_lower_in(2,33),
			in1                => s_in1(2,33),
			in2                => s_in2(2,33),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(33)
		);
	s_in1(2,33)            <= s_out1(3,33);
	s_in2(2,33)            <= s_out2(3,34);
	s_locks_lower_in(2,33) <= s_locks_lower_out(3,33);

		normal_cell_2_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,34),
			fetch              => s_fetch(2,34),
			data_in            => s_data_in(2,34),
			data_out           => s_data_out(2,34),
			out1               => s_out1(2,34),
			out2               => s_out2(2,34),
			lock_lower_row_out => s_locks_lower_out(2,34),
			lock_lower_row_in  => s_locks_lower_in(2,34),
			in1                => s_in1(2,34),
			in2                => s_in2(2,34),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(34)
		);
	s_in1(2,34)            <= s_out1(3,34);
	s_in2(2,34)            <= s_out2(3,35);
	s_locks_lower_in(2,34) <= s_locks_lower_out(3,34);

		normal_cell_2_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,35),
			fetch              => s_fetch(2,35),
			data_in            => s_data_in(2,35),
			data_out           => s_data_out(2,35),
			out1               => s_out1(2,35),
			out2               => s_out2(2,35),
			lock_lower_row_out => s_locks_lower_out(2,35),
			lock_lower_row_in  => s_locks_lower_in(2,35),
			in1                => s_in1(2,35),
			in2                => s_in2(2,35),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(35)
		);
	s_in1(2,35)            <= s_out1(3,35);
	s_in2(2,35)            <= s_out2(3,36);
	s_locks_lower_in(2,35) <= s_locks_lower_out(3,35);

		normal_cell_2_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,36),
			fetch              => s_fetch(2,36),
			data_in            => s_data_in(2,36),
			data_out           => s_data_out(2,36),
			out1               => s_out1(2,36),
			out2               => s_out2(2,36),
			lock_lower_row_out => s_locks_lower_out(2,36),
			lock_lower_row_in  => s_locks_lower_in(2,36),
			in1                => s_in1(2,36),
			in2                => s_in2(2,36),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(36)
		);
	s_in1(2,36)            <= s_out1(3,36);
	s_in2(2,36)            <= s_out2(3,37);
	s_locks_lower_in(2,36) <= s_locks_lower_out(3,36);

		normal_cell_2_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,37),
			fetch              => s_fetch(2,37),
			data_in            => s_data_in(2,37),
			data_out           => s_data_out(2,37),
			out1               => s_out1(2,37),
			out2               => s_out2(2,37),
			lock_lower_row_out => s_locks_lower_out(2,37),
			lock_lower_row_in  => s_locks_lower_in(2,37),
			in1                => s_in1(2,37),
			in2                => s_in2(2,37),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(37)
		);
	s_in1(2,37)            <= s_out1(3,37);
	s_in2(2,37)            <= s_out2(3,38);
	s_locks_lower_in(2,37) <= s_locks_lower_out(3,37);

		normal_cell_2_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,38),
			fetch              => s_fetch(2,38),
			data_in            => s_data_in(2,38),
			data_out           => s_data_out(2,38),
			out1               => s_out1(2,38),
			out2               => s_out2(2,38),
			lock_lower_row_out => s_locks_lower_out(2,38),
			lock_lower_row_in  => s_locks_lower_in(2,38),
			in1                => s_in1(2,38),
			in2                => s_in2(2,38),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(38)
		);
	s_in1(2,38)            <= s_out1(3,38);
	s_in2(2,38)            <= s_out2(3,39);
	s_locks_lower_in(2,38) <= s_locks_lower_out(3,38);

		normal_cell_2_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,39),
			fetch              => s_fetch(2,39),
			data_in            => s_data_in(2,39),
			data_out           => s_data_out(2,39),
			out1               => s_out1(2,39),
			out2               => s_out2(2,39),
			lock_lower_row_out => s_locks_lower_out(2,39),
			lock_lower_row_in  => s_locks_lower_in(2,39),
			in1                => s_in1(2,39),
			in2                => s_in2(2,39),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(39)
		);
	s_in1(2,39)            <= s_out1(3,39);
	s_in2(2,39)            <= s_out2(3,40);
	s_locks_lower_in(2,39) <= s_locks_lower_out(3,39);

		normal_cell_2_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,40),
			fetch              => s_fetch(2,40),
			data_in            => s_data_in(2,40),
			data_out           => s_data_out(2,40),
			out1               => s_out1(2,40),
			out2               => s_out2(2,40),
			lock_lower_row_out => s_locks_lower_out(2,40),
			lock_lower_row_in  => s_locks_lower_in(2,40),
			in1                => s_in1(2,40),
			in2                => s_in2(2,40),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(40)
		);
	s_in1(2,40)            <= s_out1(3,40);
	s_in2(2,40)            <= s_out2(3,41);
	s_locks_lower_in(2,40) <= s_locks_lower_out(3,40);

		normal_cell_2_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,41),
			fetch              => s_fetch(2,41),
			data_in            => s_data_in(2,41),
			data_out           => s_data_out(2,41),
			out1               => s_out1(2,41),
			out2               => s_out2(2,41),
			lock_lower_row_out => s_locks_lower_out(2,41),
			lock_lower_row_in  => s_locks_lower_in(2,41),
			in1                => s_in1(2,41),
			in2                => s_in2(2,41),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(41)
		);
	s_in1(2,41)            <= s_out1(3,41);
	s_in2(2,41)            <= s_out2(3,42);
	s_locks_lower_in(2,41) <= s_locks_lower_out(3,41);

		normal_cell_2_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,42),
			fetch              => s_fetch(2,42),
			data_in            => s_data_in(2,42),
			data_out           => s_data_out(2,42),
			out1               => s_out1(2,42),
			out2               => s_out2(2,42),
			lock_lower_row_out => s_locks_lower_out(2,42),
			lock_lower_row_in  => s_locks_lower_in(2,42),
			in1                => s_in1(2,42),
			in2                => s_in2(2,42),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(42)
		);
	s_in1(2,42)            <= s_out1(3,42);
	s_in2(2,42)            <= s_out2(3,43);
	s_locks_lower_in(2,42) <= s_locks_lower_out(3,42);

		normal_cell_2_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,43),
			fetch              => s_fetch(2,43),
			data_in            => s_data_in(2,43),
			data_out           => s_data_out(2,43),
			out1               => s_out1(2,43),
			out2               => s_out2(2,43),
			lock_lower_row_out => s_locks_lower_out(2,43),
			lock_lower_row_in  => s_locks_lower_in(2,43),
			in1                => s_in1(2,43),
			in2                => s_in2(2,43),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(43)
		);
	s_in1(2,43)            <= s_out1(3,43);
	s_in2(2,43)            <= s_out2(3,44);
	s_locks_lower_in(2,43) <= s_locks_lower_out(3,43);

		normal_cell_2_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,44),
			fetch              => s_fetch(2,44),
			data_in            => s_data_in(2,44),
			data_out           => s_data_out(2,44),
			out1               => s_out1(2,44),
			out2               => s_out2(2,44),
			lock_lower_row_out => s_locks_lower_out(2,44),
			lock_lower_row_in  => s_locks_lower_in(2,44),
			in1                => s_in1(2,44),
			in2                => s_in2(2,44),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(44)
		);
	s_in1(2,44)            <= s_out1(3,44);
	s_in2(2,44)            <= s_out2(3,45);
	s_locks_lower_in(2,44) <= s_locks_lower_out(3,44);

		normal_cell_2_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,45),
			fetch              => s_fetch(2,45),
			data_in            => s_data_in(2,45),
			data_out           => s_data_out(2,45),
			out1               => s_out1(2,45),
			out2               => s_out2(2,45),
			lock_lower_row_out => s_locks_lower_out(2,45),
			lock_lower_row_in  => s_locks_lower_in(2,45),
			in1                => s_in1(2,45),
			in2                => s_in2(2,45),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(45)
		);
	s_in1(2,45)            <= s_out1(3,45);
	s_in2(2,45)            <= s_out2(3,46);
	s_locks_lower_in(2,45) <= s_locks_lower_out(3,45);

		normal_cell_2_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,46),
			fetch              => s_fetch(2,46),
			data_in            => s_data_in(2,46),
			data_out           => s_data_out(2,46),
			out1               => s_out1(2,46),
			out2               => s_out2(2,46),
			lock_lower_row_out => s_locks_lower_out(2,46),
			lock_lower_row_in  => s_locks_lower_in(2,46),
			in1                => s_in1(2,46),
			in2                => s_in2(2,46),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(46)
		);
	s_in1(2,46)            <= s_out1(3,46);
	s_in2(2,46)            <= s_out2(3,47);
	s_locks_lower_in(2,46) <= s_locks_lower_out(3,46);

		normal_cell_2_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,47),
			fetch              => s_fetch(2,47),
			data_in            => s_data_in(2,47),
			data_out           => s_data_out(2,47),
			out1               => s_out1(2,47),
			out2               => s_out2(2,47),
			lock_lower_row_out => s_locks_lower_out(2,47),
			lock_lower_row_in  => s_locks_lower_in(2,47),
			in1                => s_in1(2,47),
			in2                => s_in2(2,47),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(47)
		);
	s_in1(2,47)            <= s_out1(3,47);
	s_in2(2,47)            <= s_out2(3,48);
	s_locks_lower_in(2,47) <= s_locks_lower_out(3,47);

		normal_cell_2_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,48),
			fetch              => s_fetch(2,48),
			data_in            => s_data_in(2,48),
			data_out           => s_data_out(2,48),
			out1               => s_out1(2,48),
			out2               => s_out2(2,48),
			lock_lower_row_out => s_locks_lower_out(2,48),
			lock_lower_row_in  => s_locks_lower_in(2,48),
			in1                => s_in1(2,48),
			in2                => s_in2(2,48),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(48)
		);
	s_in1(2,48)            <= s_out1(3,48);
	s_in2(2,48)            <= s_out2(3,49);
	s_locks_lower_in(2,48) <= s_locks_lower_out(3,48);

		normal_cell_2_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,49),
			fetch              => s_fetch(2,49),
			data_in            => s_data_in(2,49),
			data_out           => s_data_out(2,49),
			out1               => s_out1(2,49),
			out2               => s_out2(2,49),
			lock_lower_row_out => s_locks_lower_out(2,49),
			lock_lower_row_in  => s_locks_lower_in(2,49),
			in1                => s_in1(2,49),
			in2                => s_in2(2,49),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(49)
		);
	s_in1(2,49)            <= s_out1(3,49);
	s_in2(2,49)            <= s_out2(3,50);
	s_locks_lower_in(2,49) <= s_locks_lower_out(3,49);

		normal_cell_2_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,50),
			fetch              => s_fetch(2,50),
			data_in            => s_data_in(2,50),
			data_out           => s_data_out(2,50),
			out1               => s_out1(2,50),
			out2               => s_out2(2,50),
			lock_lower_row_out => s_locks_lower_out(2,50),
			lock_lower_row_in  => s_locks_lower_in(2,50),
			in1                => s_in1(2,50),
			in2                => s_in2(2,50),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(50)
		);
	s_in1(2,50)            <= s_out1(3,50);
	s_in2(2,50)            <= s_out2(3,51);
	s_locks_lower_in(2,50) <= s_locks_lower_out(3,50);

		normal_cell_2_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,51),
			fetch              => s_fetch(2,51),
			data_in            => s_data_in(2,51),
			data_out           => s_data_out(2,51),
			out1               => s_out1(2,51),
			out2               => s_out2(2,51),
			lock_lower_row_out => s_locks_lower_out(2,51),
			lock_lower_row_in  => s_locks_lower_in(2,51),
			in1                => s_in1(2,51),
			in2                => s_in2(2,51),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(51)
		);
	s_in1(2,51)            <= s_out1(3,51);
	s_in2(2,51)            <= s_out2(3,52);
	s_locks_lower_in(2,51) <= s_locks_lower_out(3,51);

		normal_cell_2_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,52),
			fetch              => s_fetch(2,52),
			data_in            => s_data_in(2,52),
			data_out           => s_data_out(2,52),
			out1               => s_out1(2,52),
			out2               => s_out2(2,52),
			lock_lower_row_out => s_locks_lower_out(2,52),
			lock_lower_row_in  => s_locks_lower_in(2,52),
			in1                => s_in1(2,52),
			in2                => s_in2(2,52),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(52)
		);
	s_in1(2,52)            <= s_out1(3,52);
	s_in2(2,52)            <= s_out2(3,53);
	s_locks_lower_in(2,52) <= s_locks_lower_out(3,52);

		normal_cell_2_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,53),
			fetch              => s_fetch(2,53),
			data_in            => s_data_in(2,53),
			data_out           => s_data_out(2,53),
			out1               => s_out1(2,53),
			out2               => s_out2(2,53),
			lock_lower_row_out => s_locks_lower_out(2,53),
			lock_lower_row_in  => s_locks_lower_in(2,53),
			in1                => s_in1(2,53),
			in2                => s_in2(2,53),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(53)
		);
	s_in1(2,53)            <= s_out1(3,53);
	s_in2(2,53)            <= s_out2(3,54);
	s_locks_lower_in(2,53) <= s_locks_lower_out(3,53);

		normal_cell_2_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,54),
			fetch              => s_fetch(2,54),
			data_in            => s_data_in(2,54),
			data_out           => s_data_out(2,54),
			out1               => s_out1(2,54),
			out2               => s_out2(2,54),
			lock_lower_row_out => s_locks_lower_out(2,54),
			lock_lower_row_in  => s_locks_lower_in(2,54),
			in1                => s_in1(2,54),
			in2                => s_in2(2,54),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(54)
		);
	s_in1(2,54)            <= s_out1(3,54);
	s_in2(2,54)            <= s_out2(3,55);
	s_locks_lower_in(2,54) <= s_locks_lower_out(3,54);

		normal_cell_2_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,55),
			fetch              => s_fetch(2,55),
			data_in            => s_data_in(2,55),
			data_out           => s_data_out(2,55),
			out1               => s_out1(2,55),
			out2               => s_out2(2,55),
			lock_lower_row_out => s_locks_lower_out(2,55),
			lock_lower_row_in  => s_locks_lower_in(2,55),
			in1                => s_in1(2,55),
			in2                => s_in2(2,55),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(55)
		);
	s_in1(2,55)            <= s_out1(3,55);
	s_in2(2,55)            <= s_out2(3,56);
	s_locks_lower_in(2,55) <= s_locks_lower_out(3,55);

		normal_cell_2_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,56),
			fetch              => s_fetch(2,56),
			data_in            => s_data_in(2,56),
			data_out           => s_data_out(2,56),
			out1               => s_out1(2,56),
			out2               => s_out2(2,56),
			lock_lower_row_out => s_locks_lower_out(2,56),
			lock_lower_row_in  => s_locks_lower_in(2,56),
			in1                => s_in1(2,56),
			in2                => s_in2(2,56),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(56)
		);
	s_in1(2,56)            <= s_out1(3,56);
	s_in2(2,56)            <= s_out2(3,57);
	s_locks_lower_in(2,56) <= s_locks_lower_out(3,56);

		normal_cell_2_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,57),
			fetch              => s_fetch(2,57),
			data_in            => s_data_in(2,57),
			data_out           => s_data_out(2,57),
			out1               => s_out1(2,57),
			out2               => s_out2(2,57),
			lock_lower_row_out => s_locks_lower_out(2,57),
			lock_lower_row_in  => s_locks_lower_in(2,57),
			in1                => s_in1(2,57),
			in2                => s_in2(2,57),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(57)
		);
	s_in1(2,57)            <= s_out1(3,57);
	s_in2(2,57)            <= s_out2(3,58);
	s_locks_lower_in(2,57) <= s_locks_lower_out(3,57);

		normal_cell_2_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,58),
			fetch              => s_fetch(2,58),
			data_in            => s_data_in(2,58),
			data_out           => s_data_out(2,58),
			out1               => s_out1(2,58),
			out2               => s_out2(2,58),
			lock_lower_row_out => s_locks_lower_out(2,58),
			lock_lower_row_in  => s_locks_lower_in(2,58),
			in1                => s_in1(2,58),
			in2                => s_in2(2,58),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(58)
		);
	s_in1(2,58)            <= s_out1(3,58);
	s_in2(2,58)            <= s_out2(3,59);
	s_locks_lower_in(2,58) <= s_locks_lower_out(3,58);

		normal_cell_2_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,59),
			fetch              => s_fetch(2,59),
			data_in            => s_data_in(2,59),
			data_out           => s_data_out(2,59),
			out1               => s_out1(2,59),
			out2               => s_out2(2,59),
			lock_lower_row_out => s_locks_lower_out(2,59),
			lock_lower_row_in  => s_locks_lower_in(2,59),
			in1                => s_in1(2,59),
			in2                => s_in2(2,59),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(59)
		);
	s_in1(2,59)            <= s_out1(3,59);
	s_in2(2,59)            <= s_out2(3,60);
	s_locks_lower_in(2,59) <= s_locks_lower_out(3,59);

		last_col_cell_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(2,60),
			fetch              => s_fetch(2,60),
			data_in            => s_data_in(2,60),
			data_out           => s_data_out(2,60),
			out1               => s_out1(2,60),
			out2               => s_out2(2,60),
			lock_lower_row_out => s_locks_lower_out(2,60),
			lock_lower_row_in  => s_locks_lower_in(2,60),
			in1                => s_in1(2,60),
			in2                => (others => '0'),
			lock_row           => s_locks(2),
			piv_found          => s_piv_found,
			row_data           => s_row_data(2),
			col_data           => s_col_data(60)
		);
	s_in1(2,60)            <= s_out1(3,60);
	s_locks_lower_in(2,60) <= s_locks_lower_out(3,60);

		normal_cell_3_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,1),
			fetch              => s_fetch(3,1),
			data_in            => s_data_in(3,1),
			data_out           => s_data_out(3,1),
			out1               => s_out1(3,1),
			out2               => s_out2(3,1),
			lock_lower_row_out => s_locks_lower_out(3,1),
			lock_lower_row_in  => s_locks_lower_in(3,1),
			in1                => s_in1(3,1),
			in2                => s_in2(3,1),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(1)
		);
	s_in1(3,1)            <= s_out1(4,1);
	s_in2(3,1)            <= s_out2(4,2);
	s_locks_lower_in(3,1) <= s_locks_lower_out(4,1);

		normal_cell_3_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,2),
			fetch              => s_fetch(3,2),
			data_in            => s_data_in(3,2),
			data_out           => s_data_out(3,2),
			out1               => s_out1(3,2),
			out2               => s_out2(3,2),
			lock_lower_row_out => s_locks_lower_out(3,2),
			lock_lower_row_in  => s_locks_lower_in(3,2),
			in1                => s_in1(3,2),
			in2                => s_in2(3,2),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(2)
		);
	s_in1(3,2)            <= s_out1(4,2);
	s_in2(3,2)            <= s_out2(4,3);
	s_locks_lower_in(3,2) <= s_locks_lower_out(4,2);

		normal_cell_3_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,3),
			fetch              => s_fetch(3,3),
			data_in            => s_data_in(3,3),
			data_out           => s_data_out(3,3),
			out1               => s_out1(3,3),
			out2               => s_out2(3,3),
			lock_lower_row_out => s_locks_lower_out(3,3),
			lock_lower_row_in  => s_locks_lower_in(3,3),
			in1                => s_in1(3,3),
			in2                => s_in2(3,3),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(3)
		);
	s_in1(3,3)            <= s_out1(4,3);
	s_in2(3,3)            <= s_out2(4,4);
	s_locks_lower_in(3,3) <= s_locks_lower_out(4,3);

		normal_cell_3_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,4),
			fetch              => s_fetch(3,4),
			data_in            => s_data_in(3,4),
			data_out           => s_data_out(3,4),
			out1               => s_out1(3,4),
			out2               => s_out2(3,4),
			lock_lower_row_out => s_locks_lower_out(3,4),
			lock_lower_row_in  => s_locks_lower_in(3,4),
			in1                => s_in1(3,4),
			in2                => s_in2(3,4),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(4)
		);
	s_in1(3,4)            <= s_out1(4,4);
	s_in2(3,4)            <= s_out2(4,5);
	s_locks_lower_in(3,4) <= s_locks_lower_out(4,4);

		normal_cell_3_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,5),
			fetch              => s_fetch(3,5),
			data_in            => s_data_in(3,5),
			data_out           => s_data_out(3,5),
			out1               => s_out1(3,5),
			out2               => s_out2(3,5),
			lock_lower_row_out => s_locks_lower_out(3,5),
			lock_lower_row_in  => s_locks_lower_in(3,5),
			in1                => s_in1(3,5),
			in2                => s_in2(3,5),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(5)
		);
	s_in1(3,5)            <= s_out1(4,5);
	s_in2(3,5)            <= s_out2(4,6);
	s_locks_lower_in(3,5) <= s_locks_lower_out(4,5);

		normal_cell_3_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,6),
			fetch              => s_fetch(3,6),
			data_in            => s_data_in(3,6),
			data_out           => s_data_out(3,6),
			out1               => s_out1(3,6),
			out2               => s_out2(3,6),
			lock_lower_row_out => s_locks_lower_out(3,6),
			lock_lower_row_in  => s_locks_lower_in(3,6),
			in1                => s_in1(3,6),
			in2                => s_in2(3,6),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(6)
		);
	s_in1(3,6)            <= s_out1(4,6);
	s_in2(3,6)            <= s_out2(4,7);
	s_locks_lower_in(3,6) <= s_locks_lower_out(4,6);

		normal_cell_3_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,7),
			fetch              => s_fetch(3,7),
			data_in            => s_data_in(3,7),
			data_out           => s_data_out(3,7),
			out1               => s_out1(3,7),
			out2               => s_out2(3,7),
			lock_lower_row_out => s_locks_lower_out(3,7),
			lock_lower_row_in  => s_locks_lower_in(3,7),
			in1                => s_in1(3,7),
			in2                => s_in2(3,7),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(7)
		);
	s_in1(3,7)            <= s_out1(4,7);
	s_in2(3,7)            <= s_out2(4,8);
	s_locks_lower_in(3,7) <= s_locks_lower_out(4,7);

		normal_cell_3_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,8),
			fetch              => s_fetch(3,8),
			data_in            => s_data_in(3,8),
			data_out           => s_data_out(3,8),
			out1               => s_out1(3,8),
			out2               => s_out2(3,8),
			lock_lower_row_out => s_locks_lower_out(3,8),
			lock_lower_row_in  => s_locks_lower_in(3,8),
			in1                => s_in1(3,8),
			in2                => s_in2(3,8),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(8)
		);
	s_in1(3,8)            <= s_out1(4,8);
	s_in2(3,8)            <= s_out2(4,9);
	s_locks_lower_in(3,8) <= s_locks_lower_out(4,8);

		normal_cell_3_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,9),
			fetch              => s_fetch(3,9),
			data_in            => s_data_in(3,9),
			data_out           => s_data_out(3,9),
			out1               => s_out1(3,9),
			out2               => s_out2(3,9),
			lock_lower_row_out => s_locks_lower_out(3,9),
			lock_lower_row_in  => s_locks_lower_in(3,9),
			in1                => s_in1(3,9),
			in2                => s_in2(3,9),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(9)
		);
	s_in1(3,9)            <= s_out1(4,9);
	s_in2(3,9)            <= s_out2(4,10);
	s_locks_lower_in(3,9) <= s_locks_lower_out(4,9);

		normal_cell_3_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,10),
			fetch              => s_fetch(3,10),
			data_in            => s_data_in(3,10),
			data_out           => s_data_out(3,10),
			out1               => s_out1(3,10),
			out2               => s_out2(3,10),
			lock_lower_row_out => s_locks_lower_out(3,10),
			lock_lower_row_in  => s_locks_lower_in(3,10),
			in1                => s_in1(3,10),
			in2                => s_in2(3,10),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(10)
		);
	s_in1(3,10)            <= s_out1(4,10);
	s_in2(3,10)            <= s_out2(4,11);
	s_locks_lower_in(3,10) <= s_locks_lower_out(4,10);

		normal_cell_3_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,11),
			fetch              => s_fetch(3,11),
			data_in            => s_data_in(3,11),
			data_out           => s_data_out(3,11),
			out1               => s_out1(3,11),
			out2               => s_out2(3,11),
			lock_lower_row_out => s_locks_lower_out(3,11),
			lock_lower_row_in  => s_locks_lower_in(3,11),
			in1                => s_in1(3,11),
			in2                => s_in2(3,11),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(11)
		);
	s_in1(3,11)            <= s_out1(4,11);
	s_in2(3,11)            <= s_out2(4,12);
	s_locks_lower_in(3,11) <= s_locks_lower_out(4,11);

		normal_cell_3_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,12),
			fetch              => s_fetch(3,12),
			data_in            => s_data_in(3,12),
			data_out           => s_data_out(3,12),
			out1               => s_out1(3,12),
			out2               => s_out2(3,12),
			lock_lower_row_out => s_locks_lower_out(3,12),
			lock_lower_row_in  => s_locks_lower_in(3,12),
			in1                => s_in1(3,12),
			in2                => s_in2(3,12),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(12)
		);
	s_in1(3,12)            <= s_out1(4,12);
	s_in2(3,12)            <= s_out2(4,13);
	s_locks_lower_in(3,12) <= s_locks_lower_out(4,12);

		normal_cell_3_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,13),
			fetch              => s_fetch(3,13),
			data_in            => s_data_in(3,13),
			data_out           => s_data_out(3,13),
			out1               => s_out1(3,13),
			out2               => s_out2(3,13),
			lock_lower_row_out => s_locks_lower_out(3,13),
			lock_lower_row_in  => s_locks_lower_in(3,13),
			in1                => s_in1(3,13),
			in2                => s_in2(3,13),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(13)
		);
	s_in1(3,13)            <= s_out1(4,13);
	s_in2(3,13)            <= s_out2(4,14);
	s_locks_lower_in(3,13) <= s_locks_lower_out(4,13);

		normal_cell_3_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,14),
			fetch              => s_fetch(3,14),
			data_in            => s_data_in(3,14),
			data_out           => s_data_out(3,14),
			out1               => s_out1(3,14),
			out2               => s_out2(3,14),
			lock_lower_row_out => s_locks_lower_out(3,14),
			lock_lower_row_in  => s_locks_lower_in(3,14),
			in1                => s_in1(3,14),
			in2                => s_in2(3,14),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(14)
		);
	s_in1(3,14)            <= s_out1(4,14);
	s_in2(3,14)            <= s_out2(4,15);
	s_locks_lower_in(3,14) <= s_locks_lower_out(4,14);

		normal_cell_3_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,15),
			fetch              => s_fetch(3,15),
			data_in            => s_data_in(3,15),
			data_out           => s_data_out(3,15),
			out1               => s_out1(3,15),
			out2               => s_out2(3,15),
			lock_lower_row_out => s_locks_lower_out(3,15),
			lock_lower_row_in  => s_locks_lower_in(3,15),
			in1                => s_in1(3,15),
			in2                => s_in2(3,15),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(15)
		);
	s_in1(3,15)            <= s_out1(4,15);
	s_in2(3,15)            <= s_out2(4,16);
	s_locks_lower_in(3,15) <= s_locks_lower_out(4,15);

		normal_cell_3_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,16),
			fetch              => s_fetch(3,16),
			data_in            => s_data_in(3,16),
			data_out           => s_data_out(3,16),
			out1               => s_out1(3,16),
			out2               => s_out2(3,16),
			lock_lower_row_out => s_locks_lower_out(3,16),
			lock_lower_row_in  => s_locks_lower_in(3,16),
			in1                => s_in1(3,16),
			in2                => s_in2(3,16),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(16)
		);
	s_in1(3,16)            <= s_out1(4,16);
	s_in2(3,16)            <= s_out2(4,17);
	s_locks_lower_in(3,16) <= s_locks_lower_out(4,16);

		normal_cell_3_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,17),
			fetch              => s_fetch(3,17),
			data_in            => s_data_in(3,17),
			data_out           => s_data_out(3,17),
			out1               => s_out1(3,17),
			out2               => s_out2(3,17),
			lock_lower_row_out => s_locks_lower_out(3,17),
			lock_lower_row_in  => s_locks_lower_in(3,17),
			in1                => s_in1(3,17),
			in2                => s_in2(3,17),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(17)
		);
	s_in1(3,17)            <= s_out1(4,17);
	s_in2(3,17)            <= s_out2(4,18);
	s_locks_lower_in(3,17) <= s_locks_lower_out(4,17);

		normal_cell_3_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,18),
			fetch              => s_fetch(3,18),
			data_in            => s_data_in(3,18),
			data_out           => s_data_out(3,18),
			out1               => s_out1(3,18),
			out2               => s_out2(3,18),
			lock_lower_row_out => s_locks_lower_out(3,18),
			lock_lower_row_in  => s_locks_lower_in(3,18),
			in1                => s_in1(3,18),
			in2                => s_in2(3,18),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(18)
		);
	s_in1(3,18)            <= s_out1(4,18);
	s_in2(3,18)            <= s_out2(4,19);
	s_locks_lower_in(3,18) <= s_locks_lower_out(4,18);

		normal_cell_3_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,19),
			fetch              => s_fetch(3,19),
			data_in            => s_data_in(3,19),
			data_out           => s_data_out(3,19),
			out1               => s_out1(3,19),
			out2               => s_out2(3,19),
			lock_lower_row_out => s_locks_lower_out(3,19),
			lock_lower_row_in  => s_locks_lower_in(3,19),
			in1                => s_in1(3,19),
			in2                => s_in2(3,19),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(19)
		);
	s_in1(3,19)            <= s_out1(4,19);
	s_in2(3,19)            <= s_out2(4,20);
	s_locks_lower_in(3,19) <= s_locks_lower_out(4,19);

		normal_cell_3_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,20),
			fetch              => s_fetch(3,20),
			data_in            => s_data_in(3,20),
			data_out           => s_data_out(3,20),
			out1               => s_out1(3,20),
			out2               => s_out2(3,20),
			lock_lower_row_out => s_locks_lower_out(3,20),
			lock_lower_row_in  => s_locks_lower_in(3,20),
			in1                => s_in1(3,20),
			in2                => s_in2(3,20),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(20)
		);
	s_in1(3,20)            <= s_out1(4,20);
	s_in2(3,20)            <= s_out2(4,21);
	s_locks_lower_in(3,20) <= s_locks_lower_out(4,20);

		normal_cell_3_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,21),
			fetch              => s_fetch(3,21),
			data_in            => s_data_in(3,21),
			data_out           => s_data_out(3,21),
			out1               => s_out1(3,21),
			out2               => s_out2(3,21),
			lock_lower_row_out => s_locks_lower_out(3,21),
			lock_lower_row_in  => s_locks_lower_in(3,21),
			in1                => s_in1(3,21),
			in2                => s_in2(3,21),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(21)
		);
	s_in1(3,21)            <= s_out1(4,21);
	s_in2(3,21)            <= s_out2(4,22);
	s_locks_lower_in(3,21) <= s_locks_lower_out(4,21);

		normal_cell_3_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,22),
			fetch              => s_fetch(3,22),
			data_in            => s_data_in(3,22),
			data_out           => s_data_out(3,22),
			out1               => s_out1(3,22),
			out2               => s_out2(3,22),
			lock_lower_row_out => s_locks_lower_out(3,22),
			lock_lower_row_in  => s_locks_lower_in(3,22),
			in1                => s_in1(3,22),
			in2                => s_in2(3,22),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(22)
		);
	s_in1(3,22)            <= s_out1(4,22);
	s_in2(3,22)            <= s_out2(4,23);
	s_locks_lower_in(3,22) <= s_locks_lower_out(4,22);

		normal_cell_3_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,23),
			fetch              => s_fetch(3,23),
			data_in            => s_data_in(3,23),
			data_out           => s_data_out(3,23),
			out1               => s_out1(3,23),
			out2               => s_out2(3,23),
			lock_lower_row_out => s_locks_lower_out(3,23),
			lock_lower_row_in  => s_locks_lower_in(3,23),
			in1                => s_in1(3,23),
			in2                => s_in2(3,23),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(23)
		);
	s_in1(3,23)            <= s_out1(4,23);
	s_in2(3,23)            <= s_out2(4,24);
	s_locks_lower_in(3,23) <= s_locks_lower_out(4,23);

		normal_cell_3_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,24),
			fetch              => s_fetch(3,24),
			data_in            => s_data_in(3,24),
			data_out           => s_data_out(3,24),
			out1               => s_out1(3,24),
			out2               => s_out2(3,24),
			lock_lower_row_out => s_locks_lower_out(3,24),
			lock_lower_row_in  => s_locks_lower_in(3,24),
			in1                => s_in1(3,24),
			in2                => s_in2(3,24),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(24)
		);
	s_in1(3,24)            <= s_out1(4,24);
	s_in2(3,24)            <= s_out2(4,25);
	s_locks_lower_in(3,24) <= s_locks_lower_out(4,24);

		normal_cell_3_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,25),
			fetch              => s_fetch(3,25),
			data_in            => s_data_in(3,25),
			data_out           => s_data_out(3,25),
			out1               => s_out1(3,25),
			out2               => s_out2(3,25),
			lock_lower_row_out => s_locks_lower_out(3,25),
			lock_lower_row_in  => s_locks_lower_in(3,25),
			in1                => s_in1(3,25),
			in2                => s_in2(3,25),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(25)
		);
	s_in1(3,25)            <= s_out1(4,25);
	s_in2(3,25)            <= s_out2(4,26);
	s_locks_lower_in(3,25) <= s_locks_lower_out(4,25);

		normal_cell_3_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,26),
			fetch              => s_fetch(3,26),
			data_in            => s_data_in(3,26),
			data_out           => s_data_out(3,26),
			out1               => s_out1(3,26),
			out2               => s_out2(3,26),
			lock_lower_row_out => s_locks_lower_out(3,26),
			lock_lower_row_in  => s_locks_lower_in(3,26),
			in1                => s_in1(3,26),
			in2                => s_in2(3,26),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(26)
		);
	s_in1(3,26)            <= s_out1(4,26);
	s_in2(3,26)            <= s_out2(4,27);
	s_locks_lower_in(3,26) <= s_locks_lower_out(4,26);

		normal_cell_3_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,27),
			fetch              => s_fetch(3,27),
			data_in            => s_data_in(3,27),
			data_out           => s_data_out(3,27),
			out1               => s_out1(3,27),
			out2               => s_out2(3,27),
			lock_lower_row_out => s_locks_lower_out(3,27),
			lock_lower_row_in  => s_locks_lower_in(3,27),
			in1                => s_in1(3,27),
			in2                => s_in2(3,27),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(27)
		);
	s_in1(3,27)            <= s_out1(4,27);
	s_in2(3,27)            <= s_out2(4,28);
	s_locks_lower_in(3,27) <= s_locks_lower_out(4,27);

		normal_cell_3_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,28),
			fetch              => s_fetch(3,28),
			data_in            => s_data_in(3,28),
			data_out           => s_data_out(3,28),
			out1               => s_out1(3,28),
			out2               => s_out2(3,28),
			lock_lower_row_out => s_locks_lower_out(3,28),
			lock_lower_row_in  => s_locks_lower_in(3,28),
			in1                => s_in1(3,28),
			in2                => s_in2(3,28),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(28)
		);
	s_in1(3,28)            <= s_out1(4,28);
	s_in2(3,28)            <= s_out2(4,29);
	s_locks_lower_in(3,28) <= s_locks_lower_out(4,28);

		normal_cell_3_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,29),
			fetch              => s_fetch(3,29),
			data_in            => s_data_in(3,29),
			data_out           => s_data_out(3,29),
			out1               => s_out1(3,29),
			out2               => s_out2(3,29),
			lock_lower_row_out => s_locks_lower_out(3,29),
			lock_lower_row_in  => s_locks_lower_in(3,29),
			in1                => s_in1(3,29),
			in2                => s_in2(3,29),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(29)
		);
	s_in1(3,29)            <= s_out1(4,29);
	s_in2(3,29)            <= s_out2(4,30);
	s_locks_lower_in(3,29) <= s_locks_lower_out(4,29);

		normal_cell_3_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,30),
			fetch              => s_fetch(3,30),
			data_in            => s_data_in(3,30),
			data_out           => s_data_out(3,30),
			out1               => s_out1(3,30),
			out2               => s_out2(3,30),
			lock_lower_row_out => s_locks_lower_out(3,30),
			lock_lower_row_in  => s_locks_lower_in(3,30),
			in1                => s_in1(3,30),
			in2                => s_in2(3,30),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(30)
		);
	s_in1(3,30)            <= s_out1(4,30);
	s_in2(3,30)            <= s_out2(4,31);
	s_locks_lower_in(3,30) <= s_locks_lower_out(4,30);

		normal_cell_3_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,31),
			fetch              => s_fetch(3,31),
			data_in            => s_data_in(3,31),
			data_out           => s_data_out(3,31),
			out1               => s_out1(3,31),
			out2               => s_out2(3,31),
			lock_lower_row_out => s_locks_lower_out(3,31),
			lock_lower_row_in  => s_locks_lower_in(3,31),
			in1                => s_in1(3,31),
			in2                => s_in2(3,31),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(31)
		);
	s_in1(3,31)            <= s_out1(4,31);
	s_in2(3,31)            <= s_out2(4,32);
	s_locks_lower_in(3,31) <= s_locks_lower_out(4,31);

		normal_cell_3_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,32),
			fetch              => s_fetch(3,32),
			data_in            => s_data_in(3,32),
			data_out           => s_data_out(3,32),
			out1               => s_out1(3,32),
			out2               => s_out2(3,32),
			lock_lower_row_out => s_locks_lower_out(3,32),
			lock_lower_row_in  => s_locks_lower_in(3,32),
			in1                => s_in1(3,32),
			in2                => s_in2(3,32),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(32)
		);
	s_in1(3,32)            <= s_out1(4,32);
	s_in2(3,32)            <= s_out2(4,33);
	s_locks_lower_in(3,32) <= s_locks_lower_out(4,32);

		normal_cell_3_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,33),
			fetch              => s_fetch(3,33),
			data_in            => s_data_in(3,33),
			data_out           => s_data_out(3,33),
			out1               => s_out1(3,33),
			out2               => s_out2(3,33),
			lock_lower_row_out => s_locks_lower_out(3,33),
			lock_lower_row_in  => s_locks_lower_in(3,33),
			in1                => s_in1(3,33),
			in2                => s_in2(3,33),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(33)
		);
	s_in1(3,33)            <= s_out1(4,33);
	s_in2(3,33)            <= s_out2(4,34);
	s_locks_lower_in(3,33) <= s_locks_lower_out(4,33);

		normal_cell_3_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,34),
			fetch              => s_fetch(3,34),
			data_in            => s_data_in(3,34),
			data_out           => s_data_out(3,34),
			out1               => s_out1(3,34),
			out2               => s_out2(3,34),
			lock_lower_row_out => s_locks_lower_out(3,34),
			lock_lower_row_in  => s_locks_lower_in(3,34),
			in1                => s_in1(3,34),
			in2                => s_in2(3,34),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(34)
		);
	s_in1(3,34)            <= s_out1(4,34);
	s_in2(3,34)            <= s_out2(4,35);
	s_locks_lower_in(3,34) <= s_locks_lower_out(4,34);

		normal_cell_3_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,35),
			fetch              => s_fetch(3,35),
			data_in            => s_data_in(3,35),
			data_out           => s_data_out(3,35),
			out1               => s_out1(3,35),
			out2               => s_out2(3,35),
			lock_lower_row_out => s_locks_lower_out(3,35),
			lock_lower_row_in  => s_locks_lower_in(3,35),
			in1                => s_in1(3,35),
			in2                => s_in2(3,35),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(35)
		);
	s_in1(3,35)            <= s_out1(4,35);
	s_in2(3,35)            <= s_out2(4,36);
	s_locks_lower_in(3,35) <= s_locks_lower_out(4,35);

		normal_cell_3_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,36),
			fetch              => s_fetch(3,36),
			data_in            => s_data_in(3,36),
			data_out           => s_data_out(3,36),
			out1               => s_out1(3,36),
			out2               => s_out2(3,36),
			lock_lower_row_out => s_locks_lower_out(3,36),
			lock_lower_row_in  => s_locks_lower_in(3,36),
			in1                => s_in1(3,36),
			in2                => s_in2(3,36),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(36)
		);
	s_in1(3,36)            <= s_out1(4,36);
	s_in2(3,36)            <= s_out2(4,37);
	s_locks_lower_in(3,36) <= s_locks_lower_out(4,36);

		normal_cell_3_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,37),
			fetch              => s_fetch(3,37),
			data_in            => s_data_in(3,37),
			data_out           => s_data_out(3,37),
			out1               => s_out1(3,37),
			out2               => s_out2(3,37),
			lock_lower_row_out => s_locks_lower_out(3,37),
			lock_lower_row_in  => s_locks_lower_in(3,37),
			in1                => s_in1(3,37),
			in2                => s_in2(3,37),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(37)
		);
	s_in1(3,37)            <= s_out1(4,37);
	s_in2(3,37)            <= s_out2(4,38);
	s_locks_lower_in(3,37) <= s_locks_lower_out(4,37);

		normal_cell_3_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,38),
			fetch              => s_fetch(3,38),
			data_in            => s_data_in(3,38),
			data_out           => s_data_out(3,38),
			out1               => s_out1(3,38),
			out2               => s_out2(3,38),
			lock_lower_row_out => s_locks_lower_out(3,38),
			lock_lower_row_in  => s_locks_lower_in(3,38),
			in1                => s_in1(3,38),
			in2                => s_in2(3,38),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(38)
		);
	s_in1(3,38)            <= s_out1(4,38);
	s_in2(3,38)            <= s_out2(4,39);
	s_locks_lower_in(3,38) <= s_locks_lower_out(4,38);

		normal_cell_3_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,39),
			fetch              => s_fetch(3,39),
			data_in            => s_data_in(3,39),
			data_out           => s_data_out(3,39),
			out1               => s_out1(3,39),
			out2               => s_out2(3,39),
			lock_lower_row_out => s_locks_lower_out(3,39),
			lock_lower_row_in  => s_locks_lower_in(3,39),
			in1                => s_in1(3,39),
			in2                => s_in2(3,39),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(39)
		);
	s_in1(3,39)            <= s_out1(4,39);
	s_in2(3,39)            <= s_out2(4,40);
	s_locks_lower_in(3,39) <= s_locks_lower_out(4,39);

		normal_cell_3_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,40),
			fetch              => s_fetch(3,40),
			data_in            => s_data_in(3,40),
			data_out           => s_data_out(3,40),
			out1               => s_out1(3,40),
			out2               => s_out2(3,40),
			lock_lower_row_out => s_locks_lower_out(3,40),
			lock_lower_row_in  => s_locks_lower_in(3,40),
			in1                => s_in1(3,40),
			in2                => s_in2(3,40),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(40)
		);
	s_in1(3,40)            <= s_out1(4,40);
	s_in2(3,40)            <= s_out2(4,41);
	s_locks_lower_in(3,40) <= s_locks_lower_out(4,40);

		normal_cell_3_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,41),
			fetch              => s_fetch(3,41),
			data_in            => s_data_in(3,41),
			data_out           => s_data_out(3,41),
			out1               => s_out1(3,41),
			out2               => s_out2(3,41),
			lock_lower_row_out => s_locks_lower_out(3,41),
			lock_lower_row_in  => s_locks_lower_in(3,41),
			in1                => s_in1(3,41),
			in2                => s_in2(3,41),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(41)
		);
	s_in1(3,41)            <= s_out1(4,41);
	s_in2(3,41)            <= s_out2(4,42);
	s_locks_lower_in(3,41) <= s_locks_lower_out(4,41);

		normal_cell_3_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,42),
			fetch              => s_fetch(3,42),
			data_in            => s_data_in(3,42),
			data_out           => s_data_out(3,42),
			out1               => s_out1(3,42),
			out2               => s_out2(3,42),
			lock_lower_row_out => s_locks_lower_out(3,42),
			lock_lower_row_in  => s_locks_lower_in(3,42),
			in1                => s_in1(3,42),
			in2                => s_in2(3,42),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(42)
		);
	s_in1(3,42)            <= s_out1(4,42);
	s_in2(3,42)            <= s_out2(4,43);
	s_locks_lower_in(3,42) <= s_locks_lower_out(4,42);

		normal_cell_3_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,43),
			fetch              => s_fetch(3,43),
			data_in            => s_data_in(3,43),
			data_out           => s_data_out(3,43),
			out1               => s_out1(3,43),
			out2               => s_out2(3,43),
			lock_lower_row_out => s_locks_lower_out(3,43),
			lock_lower_row_in  => s_locks_lower_in(3,43),
			in1                => s_in1(3,43),
			in2                => s_in2(3,43),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(43)
		);
	s_in1(3,43)            <= s_out1(4,43);
	s_in2(3,43)            <= s_out2(4,44);
	s_locks_lower_in(3,43) <= s_locks_lower_out(4,43);

		normal_cell_3_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,44),
			fetch              => s_fetch(3,44),
			data_in            => s_data_in(3,44),
			data_out           => s_data_out(3,44),
			out1               => s_out1(3,44),
			out2               => s_out2(3,44),
			lock_lower_row_out => s_locks_lower_out(3,44),
			lock_lower_row_in  => s_locks_lower_in(3,44),
			in1                => s_in1(3,44),
			in2                => s_in2(3,44),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(44)
		);
	s_in1(3,44)            <= s_out1(4,44);
	s_in2(3,44)            <= s_out2(4,45);
	s_locks_lower_in(3,44) <= s_locks_lower_out(4,44);

		normal_cell_3_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,45),
			fetch              => s_fetch(3,45),
			data_in            => s_data_in(3,45),
			data_out           => s_data_out(3,45),
			out1               => s_out1(3,45),
			out2               => s_out2(3,45),
			lock_lower_row_out => s_locks_lower_out(3,45),
			lock_lower_row_in  => s_locks_lower_in(3,45),
			in1                => s_in1(3,45),
			in2                => s_in2(3,45),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(45)
		);
	s_in1(3,45)            <= s_out1(4,45);
	s_in2(3,45)            <= s_out2(4,46);
	s_locks_lower_in(3,45) <= s_locks_lower_out(4,45);

		normal_cell_3_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,46),
			fetch              => s_fetch(3,46),
			data_in            => s_data_in(3,46),
			data_out           => s_data_out(3,46),
			out1               => s_out1(3,46),
			out2               => s_out2(3,46),
			lock_lower_row_out => s_locks_lower_out(3,46),
			lock_lower_row_in  => s_locks_lower_in(3,46),
			in1                => s_in1(3,46),
			in2                => s_in2(3,46),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(46)
		);
	s_in1(3,46)            <= s_out1(4,46);
	s_in2(3,46)            <= s_out2(4,47);
	s_locks_lower_in(3,46) <= s_locks_lower_out(4,46);

		normal_cell_3_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,47),
			fetch              => s_fetch(3,47),
			data_in            => s_data_in(3,47),
			data_out           => s_data_out(3,47),
			out1               => s_out1(3,47),
			out2               => s_out2(3,47),
			lock_lower_row_out => s_locks_lower_out(3,47),
			lock_lower_row_in  => s_locks_lower_in(3,47),
			in1                => s_in1(3,47),
			in2                => s_in2(3,47),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(47)
		);
	s_in1(3,47)            <= s_out1(4,47);
	s_in2(3,47)            <= s_out2(4,48);
	s_locks_lower_in(3,47) <= s_locks_lower_out(4,47);

		normal_cell_3_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,48),
			fetch              => s_fetch(3,48),
			data_in            => s_data_in(3,48),
			data_out           => s_data_out(3,48),
			out1               => s_out1(3,48),
			out2               => s_out2(3,48),
			lock_lower_row_out => s_locks_lower_out(3,48),
			lock_lower_row_in  => s_locks_lower_in(3,48),
			in1                => s_in1(3,48),
			in2                => s_in2(3,48),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(48)
		);
	s_in1(3,48)            <= s_out1(4,48);
	s_in2(3,48)            <= s_out2(4,49);
	s_locks_lower_in(3,48) <= s_locks_lower_out(4,48);

		normal_cell_3_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,49),
			fetch              => s_fetch(3,49),
			data_in            => s_data_in(3,49),
			data_out           => s_data_out(3,49),
			out1               => s_out1(3,49),
			out2               => s_out2(3,49),
			lock_lower_row_out => s_locks_lower_out(3,49),
			lock_lower_row_in  => s_locks_lower_in(3,49),
			in1                => s_in1(3,49),
			in2                => s_in2(3,49),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(49)
		);
	s_in1(3,49)            <= s_out1(4,49);
	s_in2(3,49)            <= s_out2(4,50);
	s_locks_lower_in(3,49) <= s_locks_lower_out(4,49);

		normal_cell_3_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,50),
			fetch              => s_fetch(3,50),
			data_in            => s_data_in(3,50),
			data_out           => s_data_out(3,50),
			out1               => s_out1(3,50),
			out2               => s_out2(3,50),
			lock_lower_row_out => s_locks_lower_out(3,50),
			lock_lower_row_in  => s_locks_lower_in(3,50),
			in1                => s_in1(3,50),
			in2                => s_in2(3,50),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(50)
		);
	s_in1(3,50)            <= s_out1(4,50);
	s_in2(3,50)            <= s_out2(4,51);
	s_locks_lower_in(3,50) <= s_locks_lower_out(4,50);

		normal_cell_3_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,51),
			fetch              => s_fetch(3,51),
			data_in            => s_data_in(3,51),
			data_out           => s_data_out(3,51),
			out1               => s_out1(3,51),
			out2               => s_out2(3,51),
			lock_lower_row_out => s_locks_lower_out(3,51),
			lock_lower_row_in  => s_locks_lower_in(3,51),
			in1                => s_in1(3,51),
			in2                => s_in2(3,51),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(51)
		);
	s_in1(3,51)            <= s_out1(4,51);
	s_in2(3,51)            <= s_out2(4,52);
	s_locks_lower_in(3,51) <= s_locks_lower_out(4,51);

		normal_cell_3_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,52),
			fetch              => s_fetch(3,52),
			data_in            => s_data_in(3,52),
			data_out           => s_data_out(3,52),
			out1               => s_out1(3,52),
			out2               => s_out2(3,52),
			lock_lower_row_out => s_locks_lower_out(3,52),
			lock_lower_row_in  => s_locks_lower_in(3,52),
			in1                => s_in1(3,52),
			in2                => s_in2(3,52),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(52)
		);
	s_in1(3,52)            <= s_out1(4,52);
	s_in2(3,52)            <= s_out2(4,53);
	s_locks_lower_in(3,52) <= s_locks_lower_out(4,52);

		normal_cell_3_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,53),
			fetch              => s_fetch(3,53),
			data_in            => s_data_in(3,53),
			data_out           => s_data_out(3,53),
			out1               => s_out1(3,53),
			out2               => s_out2(3,53),
			lock_lower_row_out => s_locks_lower_out(3,53),
			lock_lower_row_in  => s_locks_lower_in(3,53),
			in1                => s_in1(3,53),
			in2                => s_in2(3,53),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(53)
		);
	s_in1(3,53)            <= s_out1(4,53);
	s_in2(3,53)            <= s_out2(4,54);
	s_locks_lower_in(3,53) <= s_locks_lower_out(4,53);

		normal_cell_3_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,54),
			fetch              => s_fetch(3,54),
			data_in            => s_data_in(3,54),
			data_out           => s_data_out(3,54),
			out1               => s_out1(3,54),
			out2               => s_out2(3,54),
			lock_lower_row_out => s_locks_lower_out(3,54),
			lock_lower_row_in  => s_locks_lower_in(3,54),
			in1                => s_in1(3,54),
			in2                => s_in2(3,54),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(54)
		);
	s_in1(3,54)            <= s_out1(4,54);
	s_in2(3,54)            <= s_out2(4,55);
	s_locks_lower_in(3,54) <= s_locks_lower_out(4,54);

		normal_cell_3_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,55),
			fetch              => s_fetch(3,55),
			data_in            => s_data_in(3,55),
			data_out           => s_data_out(3,55),
			out1               => s_out1(3,55),
			out2               => s_out2(3,55),
			lock_lower_row_out => s_locks_lower_out(3,55),
			lock_lower_row_in  => s_locks_lower_in(3,55),
			in1                => s_in1(3,55),
			in2                => s_in2(3,55),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(55)
		);
	s_in1(3,55)            <= s_out1(4,55);
	s_in2(3,55)            <= s_out2(4,56);
	s_locks_lower_in(3,55) <= s_locks_lower_out(4,55);

		normal_cell_3_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,56),
			fetch              => s_fetch(3,56),
			data_in            => s_data_in(3,56),
			data_out           => s_data_out(3,56),
			out1               => s_out1(3,56),
			out2               => s_out2(3,56),
			lock_lower_row_out => s_locks_lower_out(3,56),
			lock_lower_row_in  => s_locks_lower_in(3,56),
			in1                => s_in1(3,56),
			in2                => s_in2(3,56),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(56)
		);
	s_in1(3,56)            <= s_out1(4,56);
	s_in2(3,56)            <= s_out2(4,57);
	s_locks_lower_in(3,56) <= s_locks_lower_out(4,56);

		normal_cell_3_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,57),
			fetch              => s_fetch(3,57),
			data_in            => s_data_in(3,57),
			data_out           => s_data_out(3,57),
			out1               => s_out1(3,57),
			out2               => s_out2(3,57),
			lock_lower_row_out => s_locks_lower_out(3,57),
			lock_lower_row_in  => s_locks_lower_in(3,57),
			in1                => s_in1(3,57),
			in2                => s_in2(3,57),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(57)
		);
	s_in1(3,57)            <= s_out1(4,57);
	s_in2(3,57)            <= s_out2(4,58);
	s_locks_lower_in(3,57) <= s_locks_lower_out(4,57);

		normal_cell_3_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,58),
			fetch              => s_fetch(3,58),
			data_in            => s_data_in(3,58),
			data_out           => s_data_out(3,58),
			out1               => s_out1(3,58),
			out2               => s_out2(3,58),
			lock_lower_row_out => s_locks_lower_out(3,58),
			lock_lower_row_in  => s_locks_lower_in(3,58),
			in1                => s_in1(3,58),
			in2                => s_in2(3,58),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(58)
		);
	s_in1(3,58)            <= s_out1(4,58);
	s_in2(3,58)            <= s_out2(4,59);
	s_locks_lower_in(3,58) <= s_locks_lower_out(4,58);

		normal_cell_3_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,59),
			fetch              => s_fetch(3,59),
			data_in            => s_data_in(3,59),
			data_out           => s_data_out(3,59),
			out1               => s_out1(3,59),
			out2               => s_out2(3,59),
			lock_lower_row_out => s_locks_lower_out(3,59),
			lock_lower_row_in  => s_locks_lower_in(3,59),
			in1                => s_in1(3,59),
			in2                => s_in2(3,59),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(59)
		);
	s_in1(3,59)            <= s_out1(4,59);
	s_in2(3,59)            <= s_out2(4,60);
	s_locks_lower_in(3,59) <= s_locks_lower_out(4,59);

		last_col_cell_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(3,60),
			fetch              => s_fetch(3,60),
			data_in            => s_data_in(3,60),
			data_out           => s_data_out(3,60),
			out1               => s_out1(3,60),
			out2               => s_out2(3,60),
			lock_lower_row_out => s_locks_lower_out(3,60),
			lock_lower_row_in  => s_locks_lower_in(3,60),
			in1                => s_in1(3,60),
			in2                => (others => '0'),
			lock_row           => s_locks(3),
			piv_found          => s_piv_found,
			row_data           => s_row_data(3),
			col_data           => s_col_data(60)
		);
	s_in1(3,60)            <= s_out1(4,60);
	s_locks_lower_in(3,60) <= s_locks_lower_out(4,60);

		normal_cell_4_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,1),
			fetch              => s_fetch(4,1),
			data_in            => s_data_in(4,1),
			data_out           => s_data_out(4,1),
			out1               => s_out1(4,1),
			out2               => s_out2(4,1),
			lock_lower_row_out => s_locks_lower_out(4,1),
			lock_lower_row_in  => s_locks_lower_in(4,1),
			in1                => s_in1(4,1),
			in2                => s_in2(4,1),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(1)
		);
	s_in1(4,1)            <= s_out1(5,1);
	s_in2(4,1)            <= s_out2(5,2);
	s_locks_lower_in(4,1) <= s_locks_lower_out(5,1);

		normal_cell_4_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,2),
			fetch              => s_fetch(4,2),
			data_in            => s_data_in(4,2),
			data_out           => s_data_out(4,2),
			out1               => s_out1(4,2),
			out2               => s_out2(4,2),
			lock_lower_row_out => s_locks_lower_out(4,2),
			lock_lower_row_in  => s_locks_lower_in(4,2),
			in1                => s_in1(4,2),
			in2                => s_in2(4,2),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(2)
		);
	s_in1(4,2)            <= s_out1(5,2);
	s_in2(4,2)            <= s_out2(5,3);
	s_locks_lower_in(4,2) <= s_locks_lower_out(5,2);

		normal_cell_4_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,3),
			fetch              => s_fetch(4,3),
			data_in            => s_data_in(4,3),
			data_out           => s_data_out(4,3),
			out1               => s_out1(4,3),
			out2               => s_out2(4,3),
			lock_lower_row_out => s_locks_lower_out(4,3),
			lock_lower_row_in  => s_locks_lower_in(4,3),
			in1                => s_in1(4,3),
			in2                => s_in2(4,3),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(3)
		);
	s_in1(4,3)            <= s_out1(5,3);
	s_in2(4,3)            <= s_out2(5,4);
	s_locks_lower_in(4,3) <= s_locks_lower_out(5,3);

		normal_cell_4_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,4),
			fetch              => s_fetch(4,4),
			data_in            => s_data_in(4,4),
			data_out           => s_data_out(4,4),
			out1               => s_out1(4,4),
			out2               => s_out2(4,4),
			lock_lower_row_out => s_locks_lower_out(4,4),
			lock_lower_row_in  => s_locks_lower_in(4,4),
			in1                => s_in1(4,4),
			in2                => s_in2(4,4),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(4)
		);
	s_in1(4,4)            <= s_out1(5,4);
	s_in2(4,4)            <= s_out2(5,5);
	s_locks_lower_in(4,4) <= s_locks_lower_out(5,4);

		normal_cell_4_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,5),
			fetch              => s_fetch(4,5),
			data_in            => s_data_in(4,5),
			data_out           => s_data_out(4,5),
			out1               => s_out1(4,5),
			out2               => s_out2(4,5),
			lock_lower_row_out => s_locks_lower_out(4,5),
			lock_lower_row_in  => s_locks_lower_in(4,5),
			in1                => s_in1(4,5),
			in2                => s_in2(4,5),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(5)
		);
	s_in1(4,5)            <= s_out1(5,5);
	s_in2(4,5)            <= s_out2(5,6);
	s_locks_lower_in(4,5) <= s_locks_lower_out(5,5);

		normal_cell_4_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,6),
			fetch              => s_fetch(4,6),
			data_in            => s_data_in(4,6),
			data_out           => s_data_out(4,6),
			out1               => s_out1(4,6),
			out2               => s_out2(4,6),
			lock_lower_row_out => s_locks_lower_out(4,6),
			lock_lower_row_in  => s_locks_lower_in(4,6),
			in1                => s_in1(4,6),
			in2                => s_in2(4,6),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(6)
		);
	s_in1(4,6)            <= s_out1(5,6);
	s_in2(4,6)            <= s_out2(5,7);
	s_locks_lower_in(4,6) <= s_locks_lower_out(5,6);

		normal_cell_4_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,7),
			fetch              => s_fetch(4,7),
			data_in            => s_data_in(4,7),
			data_out           => s_data_out(4,7),
			out1               => s_out1(4,7),
			out2               => s_out2(4,7),
			lock_lower_row_out => s_locks_lower_out(4,7),
			lock_lower_row_in  => s_locks_lower_in(4,7),
			in1                => s_in1(4,7),
			in2                => s_in2(4,7),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(7)
		);
	s_in1(4,7)            <= s_out1(5,7);
	s_in2(4,7)            <= s_out2(5,8);
	s_locks_lower_in(4,7) <= s_locks_lower_out(5,7);

		normal_cell_4_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,8),
			fetch              => s_fetch(4,8),
			data_in            => s_data_in(4,8),
			data_out           => s_data_out(4,8),
			out1               => s_out1(4,8),
			out2               => s_out2(4,8),
			lock_lower_row_out => s_locks_lower_out(4,8),
			lock_lower_row_in  => s_locks_lower_in(4,8),
			in1                => s_in1(4,8),
			in2                => s_in2(4,8),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(8)
		);
	s_in1(4,8)            <= s_out1(5,8);
	s_in2(4,8)            <= s_out2(5,9);
	s_locks_lower_in(4,8) <= s_locks_lower_out(5,8);

		normal_cell_4_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,9),
			fetch              => s_fetch(4,9),
			data_in            => s_data_in(4,9),
			data_out           => s_data_out(4,9),
			out1               => s_out1(4,9),
			out2               => s_out2(4,9),
			lock_lower_row_out => s_locks_lower_out(4,9),
			lock_lower_row_in  => s_locks_lower_in(4,9),
			in1                => s_in1(4,9),
			in2                => s_in2(4,9),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(9)
		);
	s_in1(4,9)            <= s_out1(5,9);
	s_in2(4,9)            <= s_out2(5,10);
	s_locks_lower_in(4,9) <= s_locks_lower_out(5,9);

		normal_cell_4_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,10),
			fetch              => s_fetch(4,10),
			data_in            => s_data_in(4,10),
			data_out           => s_data_out(4,10),
			out1               => s_out1(4,10),
			out2               => s_out2(4,10),
			lock_lower_row_out => s_locks_lower_out(4,10),
			lock_lower_row_in  => s_locks_lower_in(4,10),
			in1                => s_in1(4,10),
			in2                => s_in2(4,10),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(10)
		);
	s_in1(4,10)            <= s_out1(5,10);
	s_in2(4,10)            <= s_out2(5,11);
	s_locks_lower_in(4,10) <= s_locks_lower_out(5,10);

		normal_cell_4_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,11),
			fetch              => s_fetch(4,11),
			data_in            => s_data_in(4,11),
			data_out           => s_data_out(4,11),
			out1               => s_out1(4,11),
			out2               => s_out2(4,11),
			lock_lower_row_out => s_locks_lower_out(4,11),
			lock_lower_row_in  => s_locks_lower_in(4,11),
			in1                => s_in1(4,11),
			in2                => s_in2(4,11),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(11)
		);
	s_in1(4,11)            <= s_out1(5,11);
	s_in2(4,11)            <= s_out2(5,12);
	s_locks_lower_in(4,11) <= s_locks_lower_out(5,11);

		normal_cell_4_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,12),
			fetch              => s_fetch(4,12),
			data_in            => s_data_in(4,12),
			data_out           => s_data_out(4,12),
			out1               => s_out1(4,12),
			out2               => s_out2(4,12),
			lock_lower_row_out => s_locks_lower_out(4,12),
			lock_lower_row_in  => s_locks_lower_in(4,12),
			in1                => s_in1(4,12),
			in2                => s_in2(4,12),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(12)
		);
	s_in1(4,12)            <= s_out1(5,12);
	s_in2(4,12)            <= s_out2(5,13);
	s_locks_lower_in(4,12) <= s_locks_lower_out(5,12);

		normal_cell_4_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,13),
			fetch              => s_fetch(4,13),
			data_in            => s_data_in(4,13),
			data_out           => s_data_out(4,13),
			out1               => s_out1(4,13),
			out2               => s_out2(4,13),
			lock_lower_row_out => s_locks_lower_out(4,13),
			lock_lower_row_in  => s_locks_lower_in(4,13),
			in1                => s_in1(4,13),
			in2                => s_in2(4,13),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(13)
		);
	s_in1(4,13)            <= s_out1(5,13);
	s_in2(4,13)            <= s_out2(5,14);
	s_locks_lower_in(4,13) <= s_locks_lower_out(5,13);

		normal_cell_4_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,14),
			fetch              => s_fetch(4,14),
			data_in            => s_data_in(4,14),
			data_out           => s_data_out(4,14),
			out1               => s_out1(4,14),
			out2               => s_out2(4,14),
			lock_lower_row_out => s_locks_lower_out(4,14),
			lock_lower_row_in  => s_locks_lower_in(4,14),
			in1                => s_in1(4,14),
			in2                => s_in2(4,14),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(14)
		);
	s_in1(4,14)            <= s_out1(5,14);
	s_in2(4,14)            <= s_out2(5,15);
	s_locks_lower_in(4,14) <= s_locks_lower_out(5,14);

		normal_cell_4_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,15),
			fetch              => s_fetch(4,15),
			data_in            => s_data_in(4,15),
			data_out           => s_data_out(4,15),
			out1               => s_out1(4,15),
			out2               => s_out2(4,15),
			lock_lower_row_out => s_locks_lower_out(4,15),
			lock_lower_row_in  => s_locks_lower_in(4,15),
			in1                => s_in1(4,15),
			in2                => s_in2(4,15),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(15)
		);
	s_in1(4,15)            <= s_out1(5,15);
	s_in2(4,15)            <= s_out2(5,16);
	s_locks_lower_in(4,15) <= s_locks_lower_out(5,15);

		normal_cell_4_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,16),
			fetch              => s_fetch(4,16),
			data_in            => s_data_in(4,16),
			data_out           => s_data_out(4,16),
			out1               => s_out1(4,16),
			out2               => s_out2(4,16),
			lock_lower_row_out => s_locks_lower_out(4,16),
			lock_lower_row_in  => s_locks_lower_in(4,16),
			in1                => s_in1(4,16),
			in2                => s_in2(4,16),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(16)
		);
	s_in1(4,16)            <= s_out1(5,16);
	s_in2(4,16)            <= s_out2(5,17);
	s_locks_lower_in(4,16) <= s_locks_lower_out(5,16);

		normal_cell_4_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,17),
			fetch              => s_fetch(4,17),
			data_in            => s_data_in(4,17),
			data_out           => s_data_out(4,17),
			out1               => s_out1(4,17),
			out2               => s_out2(4,17),
			lock_lower_row_out => s_locks_lower_out(4,17),
			lock_lower_row_in  => s_locks_lower_in(4,17),
			in1                => s_in1(4,17),
			in2                => s_in2(4,17),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(17)
		);
	s_in1(4,17)            <= s_out1(5,17);
	s_in2(4,17)            <= s_out2(5,18);
	s_locks_lower_in(4,17) <= s_locks_lower_out(5,17);

		normal_cell_4_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,18),
			fetch              => s_fetch(4,18),
			data_in            => s_data_in(4,18),
			data_out           => s_data_out(4,18),
			out1               => s_out1(4,18),
			out2               => s_out2(4,18),
			lock_lower_row_out => s_locks_lower_out(4,18),
			lock_lower_row_in  => s_locks_lower_in(4,18),
			in1                => s_in1(4,18),
			in2                => s_in2(4,18),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(18)
		);
	s_in1(4,18)            <= s_out1(5,18);
	s_in2(4,18)            <= s_out2(5,19);
	s_locks_lower_in(4,18) <= s_locks_lower_out(5,18);

		normal_cell_4_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,19),
			fetch              => s_fetch(4,19),
			data_in            => s_data_in(4,19),
			data_out           => s_data_out(4,19),
			out1               => s_out1(4,19),
			out2               => s_out2(4,19),
			lock_lower_row_out => s_locks_lower_out(4,19),
			lock_lower_row_in  => s_locks_lower_in(4,19),
			in1                => s_in1(4,19),
			in2                => s_in2(4,19),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(19)
		);
	s_in1(4,19)            <= s_out1(5,19);
	s_in2(4,19)            <= s_out2(5,20);
	s_locks_lower_in(4,19) <= s_locks_lower_out(5,19);

		normal_cell_4_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,20),
			fetch              => s_fetch(4,20),
			data_in            => s_data_in(4,20),
			data_out           => s_data_out(4,20),
			out1               => s_out1(4,20),
			out2               => s_out2(4,20),
			lock_lower_row_out => s_locks_lower_out(4,20),
			lock_lower_row_in  => s_locks_lower_in(4,20),
			in1                => s_in1(4,20),
			in2                => s_in2(4,20),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(20)
		);
	s_in1(4,20)            <= s_out1(5,20);
	s_in2(4,20)            <= s_out2(5,21);
	s_locks_lower_in(4,20) <= s_locks_lower_out(5,20);

		normal_cell_4_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,21),
			fetch              => s_fetch(4,21),
			data_in            => s_data_in(4,21),
			data_out           => s_data_out(4,21),
			out1               => s_out1(4,21),
			out2               => s_out2(4,21),
			lock_lower_row_out => s_locks_lower_out(4,21),
			lock_lower_row_in  => s_locks_lower_in(4,21),
			in1                => s_in1(4,21),
			in2                => s_in2(4,21),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(21)
		);
	s_in1(4,21)            <= s_out1(5,21);
	s_in2(4,21)            <= s_out2(5,22);
	s_locks_lower_in(4,21) <= s_locks_lower_out(5,21);

		normal_cell_4_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,22),
			fetch              => s_fetch(4,22),
			data_in            => s_data_in(4,22),
			data_out           => s_data_out(4,22),
			out1               => s_out1(4,22),
			out2               => s_out2(4,22),
			lock_lower_row_out => s_locks_lower_out(4,22),
			lock_lower_row_in  => s_locks_lower_in(4,22),
			in1                => s_in1(4,22),
			in2                => s_in2(4,22),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(22)
		);
	s_in1(4,22)            <= s_out1(5,22);
	s_in2(4,22)            <= s_out2(5,23);
	s_locks_lower_in(4,22) <= s_locks_lower_out(5,22);

		normal_cell_4_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,23),
			fetch              => s_fetch(4,23),
			data_in            => s_data_in(4,23),
			data_out           => s_data_out(4,23),
			out1               => s_out1(4,23),
			out2               => s_out2(4,23),
			lock_lower_row_out => s_locks_lower_out(4,23),
			lock_lower_row_in  => s_locks_lower_in(4,23),
			in1                => s_in1(4,23),
			in2                => s_in2(4,23),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(23)
		);
	s_in1(4,23)            <= s_out1(5,23);
	s_in2(4,23)            <= s_out2(5,24);
	s_locks_lower_in(4,23) <= s_locks_lower_out(5,23);

		normal_cell_4_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,24),
			fetch              => s_fetch(4,24),
			data_in            => s_data_in(4,24),
			data_out           => s_data_out(4,24),
			out1               => s_out1(4,24),
			out2               => s_out2(4,24),
			lock_lower_row_out => s_locks_lower_out(4,24),
			lock_lower_row_in  => s_locks_lower_in(4,24),
			in1                => s_in1(4,24),
			in2                => s_in2(4,24),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(24)
		);
	s_in1(4,24)            <= s_out1(5,24);
	s_in2(4,24)            <= s_out2(5,25);
	s_locks_lower_in(4,24) <= s_locks_lower_out(5,24);

		normal_cell_4_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,25),
			fetch              => s_fetch(4,25),
			data_in            => s_data_in(4,25),
			data_out           => s_data_out(4,25),
			out1               => s_out1(4,25),
			out2               => s_out2(4,25),
			lock_lower_row_out => s_locks_lower_out(4,25),
			lock_lower_row_in  => s_locks_lower_in(4,25),
			in1                => s_in1(4,25),
			in2                => s_in2(4,25),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(25)
		);
	s_in1(4,25)            <= s_out1(5,25);
	s_in2(4,25)            <= s_out2(5,26);
	s_locks_lower_in(4,25) <= s_locks_lower_out(5,25);

		normal_cell_4_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,26),
			fetch              => s_fetch(4,26),
			data_in            => s_data_in(4,26),
			data_out           => s_data_out(4,26),
			out1               => s_out1(4,26),
			out2               => s_out2(4,26),
			lock_lower_row_out => s_locks_lower_out(4,26),
			lock_lower_row_in  => s_locks_lower_in(4,26),
			in1                => s_in1(4,26),
			in2                => s_in2(4,26),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(26)
		);
	s_in1(4,26)            <= s_out1(5,26);
	s_in2(4,26)            <= s_out2(5,27);
	s_locks_lower_in(4,26) <= s_locks_lower_out(5,26);

		normal_cell_4_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,27),
			fetch              => s_fetch(4,27),
			data_in            => s_data_in(4,27),
			data_out           => s_data_out(4,27),
			out1               => s_out1(4,27),
			out2               => s_out2(4,27),
			lock_lower_row_out => s_locks_lower_out(4,27),
			lock_lower_row_in  => s_locks_lower_in(4,27),
			in1                => s_in1(4,27),
			in2                => s_in2(4,27),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(27)
		);
	s_in1(4,27)            <= s_out1(5,27);
	s_in2(4,27)            <= s_out2(5,28);
	s_locks_lower_in(4,27) <= s_locks_lower_out(5,27);

		normal_cell_4_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,28),
			fetch              => s_fetch(4,28),
			data_in            => s_data_in(4,28),
			data_out           => s_data_out(4,28),
			out1               => s_out1(4,28),
			out2               => s_out2(4,28),
			lock_lower_row_out => s_locks_lower_out(4,28),
			lock_lower_row_in  => s_locks_lower_in(4,28),
			in1                => s_in1(4,28),
			in2                => s_in2(4,28),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(28)
		);
	s_in1(4,28)            <= s_out1(5,28);
	s_in2(4,28)            <= s_out2(5,29);
	s_locks_lower_in(4,28) <= s_locks_lower_out(5,28);

		normal_cell_4_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,29),
			fetch              => s_fetch(4,29),
			data_in            => s_data_in(4,29),
			data_out           => s_data_out(4,29),
			out1               => s_out1(4,29),
			out2               => s_out2(4,29),
			lock_lower_row_out => s_locks_lower_out(4,29),
			lock_lower_row_in  => s_locks_lower_in(4,29),
			in1                => s_in1(4,29),
			in2                => s_in2(4,29),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(29)
		);
	s_in1(4,29)            <= s_out1(5,29);
	s_in2(4,29)            <= s_out2(5,30);
	s_locks_lower_in(4,29) <= s_locks_lower_out(5,29);

		normal_cell_4_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,30),
			fetch              => s_fetch(4,30),
			data_in            => s_data_in(4,30),
			data_out           => s_data_out(4,30),
			out1               => s_out1(4,30),
			out2               => s_out2(4,30),
			lock_lower_row_out => s_locks_lower_out(4,30),
			lock_lower_row_in  => s_locks_lower_in(4,30),
			in1                => s_in1(4,30),
			in2                => s_in2(4,30),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(30)
		);
	s_in1(4,30)            <= s_out1(5,30);
	s_in2(4,30)            <= s_out2(5,31);
	s_locks_lower_in(4,30) <= s_locks_lower_out(5,30);

		normal_cell_4_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,31),
			fetch              => s_fetch(4,31),
			data_in            => s_data_in(4,31),
			data_out           => s_data_out(4,31),
			out1               => s_out1(4,31),
			out2               => s_out2(4,31),
			lock_lower_row_out => s_locks_lower_out(4,31),
			lock_lower_row_in  => s_locks_lower_in(4,31),
			in1                => s_in1(4,31),
			in2                => s_in2(4,31),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(31)
		);
	s_in1(4,31)            <= s_out1(5,31);
	s_in2(4,31)            <= s_out2(5,32);
	s_locks_lower_in(4,31) <= s_locks_lower_out(5,31);

		normal_cell_4_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,32),
			fetch              => s_fetch(4,32),
			data_in            => s_data_in(4,32),
			data_out           => s_data_out(4,32),
			out1               => s_out1(4,32),
			out2               => s_out2(4,32),
			lock_lower_row_out => s_locks_lower_out(4,32),
			lock_lower_row_in  => s_locks_lower_in(4,32),
			in1                => s_in1(4,32),
			in2                => s_in2(4,32),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(32)
		);
	s_in1(4,32)            <= s_out1(5,32);
	s_in2(4,32)            <= s_out2(5,33);
	s_locks_lower_in(4,32) <= s_locks_lower_out(5,32);

		normal_cell_4_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,33),
			fetch              => s_fetch(4,33),
			data_in            => s_data_in(4,33),
			data_out           => s_data_out(4,33),
			out1               => s_out1(4,33),
			out2               => s_out2(4,33),
			lock_lower_row_out => s_locks_lower_out(4,33),
			lock_lower_row_in  => s_locks_lower_in(4,33),
			in1                => s_in1(4,33),
			in2                => s_in2(4,33),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(33)
		);
	s_in1(4,33)            <= s_out1(5,33);
	s_in2(4,33)            <= s_out2(5,34);
	s_locks_lower_in(4,33) <= s_locks_lower_out(5,33);

		normal_cell_4_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,34),
			fetch              => s_fetch(4,34),
			data_in            => s_data_in(4,34),
			data_out           => s_data_out(4,34),
			out1               => s_out1(4,34),
			out2               => s_out2(4,34),
			lock_lower_row_out => s_locks_lower_out(4,34),
			lock_lower_row_in  => s_locks_lower_in(4,34),
			in1                => s_in1(4,34),
			in2                => s_in2(4,34),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(34)
		);
	s_in1(4,34)            <= s_out1(5,34);
	s_in2(4,34)            <= s_out2(5,35);
	s_locks_lower_in(4,34) <= s_locks_lower_out(5,34);

		normal_cell_4_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,35),
			fetch              => s_fetch(4,35),
			data_in            => s_data_in(4,35),
			data_out           => s_data_out(4,35),
			out1               => s_out1(4,35),
			out2               => s_out2(4,35),
			lock_lower_row_out => s_locks_lower_out(4,35),
			lock_lower_row_in  => s_locks_lower_in(4,35),
			in1                => s_in1(4,35),
			in2                => s_in2(4,35),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(35)
		);
	s_in1(4,35)            <= s_out1(5,35);
	s_in2(4,35)            <= s_out2(5,36);
	s_locks_lower_in(4,35) <= s_locks_lower_out(5,35);

		normal_cell_4_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,36),
			fetch              => s_fetch(4,36),
			data_in            => s_data_in(4,36),
			data_out           => s_data_out(4,36),
			out1               => s_out1(4,36),
			out2               => s_out2(4,36),
			lock_lower_row_out => s_locks_lower_out(4,36),
			lock_lower_row_in  => s_locks_lower_in(4,36),
			in1                => s_in1(4,36),
			in2                => s_in2(4,36),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(36)
		);
	s_in1(4,36)            <= s_out1(5,36);
	s_in2(4,36)            <= s_out2(5,37);
	s_locks_lower_in(4,36) <= s_locks_lower_out(5,36);

		normal_cell_4_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,37),
			fetch              => s_fetch(4,37),
			data_in            => s_data_in(4,37),
			data_out           => s_data_out(4,37),
			out1               => s_out1(4,37),
			out2               => s_out2(4,37),
			lock_lower_row_out => s_locks_lower_out(4,37),
			lock_lower_row_in  => s_locks_lower_in(4,37),
			in1                => s_in1(4,37),
			in2                => s_in2(4,37),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(37)
		);
	s_in1(4,37)            <= s_out1(5,37);
	s_in2(4,37)            <= s_out2(5,38);
	s_locks_lower_in(4,37) <= s_locks_lower_out(5,37);

		normal_cell_4_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,38),
			fetch              => s_fetch(4,38),
			data_in            => s_data_in(4,38),
			data_out           => s_data_out(4,38),
			out1               => s_out1(4,38),
			out2               => s_out2(4,38),
			lock_lower_row_out => s_locks_lower_out(4,38),
			lock_lower_row_in  => s_locks_lower_in(4,38),
			in1                => s_in1(4,38),
			in2                => s_in2(4,38),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(38)
		);
	s_in1(4,38)            <= s_out1(5,38);
	s_in2(4,38)            <= s_out2(5,39);
	s_locks_lower_in(4,38) <= s_locks_lower_out(5,38);

		normal_cell_4_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,39),
			fetch              => s_fetch(4,39),
			data_in            => s_data_in(4,39),
			data_out           => s_data_out(4,39),
			out1               => s_out1(4,39),
			out2               => s_out2(4,39),
			lock_lower_row_out => s_locks_lower_out(4,39),
			lock_lower_row_in  => s_locks_lower_in(4,39),
			in1                => s_in1(4,39),
			in2                => s_in2(4,39),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(39)
		);
	s_in1(4,39)            <= s_out1(5,39);
	s_in2(4,39)            <= s_out2(5,40);
	s_locks_lower_in(4,39) <= s_locks_lower_out(5,39);

		normal_cell_4_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,40),
			fetch              => s_fetch(4,40),
			data_in            => s_data_in(4,40),
			data_out           => s_data_out(4,40),
			out1               => s_out1(4,40),
			out2               => s_out2(4,40),
			lock_lower_row_out => s_locks_lower_out(4,40),
			lock_lower_row_in  => s_locks_lower_in(4,40),
			in1                => s_in1(4,40),
			in2                => s_in2(4,40),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(40)
		);
	s_in1(4,40)            <= s_out1(5,40);
	s_in2(4,40)            <= s_out2(5,41);
	s_locks_lower_in(4,40) <= s_locks_lower_out(5,40);

		normal_cell_4_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,41),
			fetch              => s_fetch(4,41),
			data_in            => s_data_in(4,41),
			data_out           => s_data_out(4,41),
			out1               => s_out1(4,41),
			out2               => s_out2(4,41),
			lock_lower_row_out => s_locks_lower_out(4,41),
			lock_lower_row_in  => s_locks_lower_in(4,41),
			in1                => s_in1(4,41),
			in2                => s_in2(4,41),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(41)
		);
	s_in1(4,41)            <= s_out1(5,41);
	s_in2(4,41)            <= s_out2(5,42);
	s_locks_lower_in(4,41) <= s_locks_lower_out(5,41);

		normal_cell_4_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,42),
			fetch              => s_fetch(4,42),
			data_in            => s_data_in(4,42),
			data_out           => s_data_out(4,42),
			out1               => s_out1(4,42),
			out2               => s_out2(4,42),
			lock_lower_row_out => s_locks_lower_out(4,42),
			lock_lower_row_in  => s_locks_lower_in(4,42),
			in1                => s_in1(4,42),
			in2                => s_in2(4,42),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(42)
		);
	s_in1(4,42)            <= s_out1(5,42);
	s_in2(4,42)            <= s_out2(5,43);
	s_locks_lower_in(4,42) <= s_locks_lower_out(5,42);

		normal_cell_4_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,43),
			fetch              => s_fetch(4,43),
			data_in            => s_data_in(4,43),
			data_out           => s_data_out(4,43),
			out1               => s_out1(4,43),
			out2               => s_out2(4,43),
			lock_lower_row_out => s_locks_lower_out(4,43),
			lock_lower_row_in  => s_locks_lower_in(4,43),
			in1                => s_in1(4,43),
			in2                => s_in2(4,43),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(43)
		);
	s_in1(4,43)            <= s_out1(5,43);
	s_in2(4,43)            <= s_out2(5,44);
	s_locks_lower_in(4,43) <= s_locks_lower_out(5,43);

		normal_cell_4_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,44),
			fetch              => s_fetch(4,44),
			data_in            => s_data_in(4,44),
			data_out           => s_data_out(4,44),
			out1               => s_out1(4,44),
			out2               => s_out2(4,44),
			lock_lower_row_out => s_locks_lower_out(4,44),
			lock_lower_row_in  => s_locks_lower_in(4,44),
			in1                => s_in1(4,44),
			in2                => s_in2(4,44),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(44)
		);
	s_in1(4,44)            <= s_out1(5,44);
	s_in2(4,44)            <= s_out2(5,45);
	s_locks_lower_in(4,44) <= s_locks_lower_out(5,44);

		normal_cell_4_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,45),
			fetch              => s_fetch(4,45),
			data_in            => s_data_in(4,45),
			data_out           => s_data_out(4,45),
			out1               => s_out1(4,45),
			out2               => s_out2(4,45),
			lock_lower_row_out => s_locks_lower_out(4,45),
			lock_lower_row_in  => s_locks_lower_in(4,45),
			in1                => s_in1(4,45),
			in2                => s_in2(4,45),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(45)
		);
	s_in1(4,45)            <= s_out1(5,45);
	s_in2(4,45)            <= s_out2(5,46);
	s_locks_lower_in(4,45) <= s_locks_lower_out(5,45);

		normal_cell_4_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,46),
			fetch              => s_fetch(4,46),
			data_in            => s_data_in(4,46),
			data_out           => s_data_out(4,46),
			out1               => s_out1(4,46),
			out2               => s_out2(4,46),
			lock_lower_row_out => s_locks_lower_out(4,46),
			lock_lower_row_in  => s_locks_lower_in(4,46),
			in1                => s_in1(4,46),
			in2                => s_in2(4,46),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(46)
		);
	s_in1(4,46)            <= s_out1(5,46);
	s_in2(4,46)            <= s_out2(5,47);
	s_locks_lower_in(4,46) <= s_locks_lower_out(5,46);

		normal_cell_4_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,47),
			fetch              => s_fetch(4,47),
			data_in            => s_data_in(4,47),
			data_out           => s_data_out(4,47),
			out1               => s_out1(4,47),
			out2               => s_out2(4,47),
			lock_lower_row_out => s_locks_lower_out(4,47),
			lock_lower_row_in  => s_locks_lower_in(4,47),
			in1                => s_in1(4,47),
			in2                => s_in2(4,47),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(47)
		);
	s_in1(4,47)            <= s_out1(5,47);
	s_in2(4,47)            <= s_out2(5,48);
	s_locks_lower_in(4,47) <= s_locks_lower_out(5,47);

		normal_cell_4_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,48),
			fetch              => s_fetch(4,48),
			data_in            => s_data_in(4,48),
			data_out           => s_data_out(4,48),
			out1               => s_out1(4,48),
			out2               => s_out2(4,48),
			lock_lower_row_out => s_locks_lower_out(4,48),
			lock_lower_row_in  => s_locks_lower_in(4,48),
			in1                => s_in1(4,48),
			in2                => s_in2(4,48),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(48)
		);
	s_in1(4,48)            <= s_out1(5,48);
	s_in2(4,48)            <= s_out2(5,49);
	s_locks_lower_in(4,48) <= s_locks_lower_out(5,48);

		normal_cell_4_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,49),
			fetch              => s_fetch(4,49),
			data_in            => s_data_in(4,49),
			data_out           => s_data_out(4,49),
			out1               => s_out1(4,49),
			out2               => s_out2(4,49),
			lock_lower_row_out => s_locks_lower_out(4,49),
			lock_lower_row_in  => s_locks_lower_in(4,49),
			in1                => s_in1(4,49),
			in2                => s_in2(4,49),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(49)
		);
	s_in1(4,49)            <= s_out1(5,49);
	s_in2(4,49)            <= s_out2(5,50);
	s_locks_lower_in(4,49) <= s_locks_lower_out(5,49);

		normal_cell_4_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,50),
			fetch              => s_fetch(4,50),
			data_in            => s_data_in(4,50),
			data_out           => s_data_out(4,50),
			out1               => s_out1(4,50),
			out2               => s_out2(4,50),
			lock_lower_row_out => s_locks_lower_out(4,50),
			lock_lower_row_in  => s_locks_lower_in(4,50),
			in1                => s_in1(4,50),
			in2                => s_in2(4,50),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(50)
		);
	s_in1(4,50)            <= s_out1(5,50);
	s_in2(4,50)            <= s_out2(5,51);
	s_locks_lower_in(4,50) <= s_locks_lower_out(5,50);

		normal_cell_4_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,51),
			fetch              => s_fetch(4,51),
			data_in            => s_data_in(4,51),
			data_out           => s_data_out(4,51),
			out1               => s_out1(4,51),
			out2               => s_out2(4,51),
			lock_lower_row_out => s_locks_lower_out(4,51),
			lock_lower_row_in  => s_locks_lower_in(4,51),
			in1                => s_in1(4,51),
			in2                => s_in2(4,51),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(51)
		);
	s_in1(4,51)            <= s_out1(5,51);
	s_in2(4,51)            <= s_out2(5,52);
	s_locks_lower_in(4,51) <= s_locks_lower_out(5,51);

		normal_cell_4_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,52),
			fetch              => s_fetch(4,52),
			data_in            => s_data_in(4,52),
			data_out           => s_data_out(4,52),
			out1               => s_out1(4,52),
			out2               => s_out2(4,52),
			lock_lower_row_out => s_locks_lower_out(4,52),
			lock_lower_row_in  => s_locks_lower_in(4,52),
			in1                => s_in1(4,52),
			in2                => s_in2(4,52),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(52)
		);
	s_in1(4,52)            <= s_out1(5,52);
	s_in2(4,52)            <= s_out2(5,53);
	s_locks_lower_in(4,52) <= s_locks_lower_out(5,52);

		normal_cell_4_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,53),
			fetch              => s_fetch(4,53),
			data_in            => s_data_in(4,53),
			data_out           => s_data_out(4,53),
			out1               => s_out1(4,53),
			out2               => s_out2(4,53),
			lock_lower_row_out => s_locks_lower_out(4,53),
			lock_lower_row_in  => s_locks_lower_in(4,53),
			in1                => s_in1(4,53),
			in2                => s_in2(4,53),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(53)
		);
	s_in1(4,53)            <= s_out1(5,53);
	s_in2(4,53)            <= s_out2(5,54);
	s_locks_lower_in(4,53) <= s_locks_lower_out(5,53);

		normal_cell_4_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,54),
			fetch              => s_fetch(4,54),
			data_in            => s_data_in(4,54),
			data_out           => s_data_out(4,54),
			out1               => s_out1(4,54),
			out2               => s_out2(4,54),
			lock_lower_row_out => s_locks_lower_out(4,54),
			lock_lower_row_in  => s_locks_lower_in(4,54),
			in1                => s_in1(4,54),
			in2                => s_in2(4,54),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(54)
		);
	s_in1(4,54)            <= s_out1(5,54);
	s_in2(4,54)            <= s_out2(5,55);
	s_locks_lower_in(4,54) <= s_locks_lower_out(5,54);

		normal_cell_4_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,55),
			fetch              => s_fetch(4,55),
			data_in            => s_data_in(4,55),
			data_out           => s_data_out(4,55),
			out1               => s_out1(4,55),
			out2               => s_out2(4,55),
			lock_lower_row_out => s_locks_lower_out(4,55),
			lock_lower_row_in  => s_locks_lower_in(4,55),
			in1                => s_in1(4,55),
			in2                => s_in2(4,55),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(55)
		);
	s_in1(4,55)            <= s_out1(5,55);
	s_in2(4,55)            <= s_out2(5,56);
	s_locks_lower_in(4,55) <= s_locks_lower_out(5,55);

		normal_cell_4_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,56),
			fetch              => s_fetch(4,56),
			data_in            => s_data_in(4,56),
			data_out           => s_data_out(4,56),
			out1               => s_out1(4,56),
			out2               => s_out2(4,56),
			lock_lower_row_out => s_locks_lower_out(4,56),
			lock_lower_row_in  => s_locks_lower_in(4,56),
			in1                => s_in1(4,56),
			in2                => s_in2(4,56),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(56)
		);
	s_in1(4,56)            <= s_out1(5,56);
	s_in2(4,56)            <= s_out2(5,57);
	s_locks_lower_in(4,56) <= s_locks_lower_out(5,56);

		normal_cell_4_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,57),
			fetch              => s_fetch(4,57),
			data_in            => s_data_in(4,57),
			data_out           => s_data_out(4,57),
			out1               => s_out1(4,57),
			out2               => s_out2(4,57),
			lock_lower_row_out => s_locks_lower_out(4,57),
			lock_lower_row_in  => s_locks_lower_in(4,57),
			in1                => s_in1(4,57),
			in2                => s_in2(4,57),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(57)
		);
	s_in1(4,57)            <= s_out1(5,57);
	s_in2(4,57)            <= s_out2(5,58);
	s_locks_lower_in(4,57) <= s_locks_lower_out(5,57);

		normal_cell_4_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,58),
			fetch              => s_fetch(4,58),
			data_in            => s_data_in(4,58),
			data_out           => s_data_out(4,58),
			out1               => s_out1(4,58),
			out2               => s_out2(4,58),
			lock_lower_row_out => s_locks_lower_out(4,58),
			lock_lower_row_in  => s_locks_lower_in(4,58),
			in1                => s_in1(4,58),
			in2                => s_in2(4,58),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(58)
		);
	s_in1(4,58)            <= s_out1(5,58);
	s_in2(4,58)            <= s_out2(5,59);
	s_locks_lower_in(4,58) <= s_locks_lower_out(5,58);

		normal_cell_4_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,59),
			fetch              => s_fetch(4,59),
			data_in            => s_data_in(4,59),
			data_out           => s_data_out(4,59),
			out1               => s_out1(4,59),
			out2               => s_out2(4,59),
			lock_lower_row_out => s_locks_lower_out(4,59),
			lock_lower_row_in  => s_locks_lower_in(4,59),
			in1                => s_in1(4,59),
			in2                => s_in2(4,59),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(59)
		);
	s_in1(4,59)            <= s_out1(5,59);
	s_in2(4,59)            <= s_out2(5,60);
	s_locks_lower_in(4,59) <= s_locks_lower_out(5,59);

		last_col_cell_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(4,60),
			fetch              => s_fetch(4,60),
			data_in            => s_data_in(4,60),
			data_out           => s_data_out(4,60),
			out1               => s_out1(4,60),
			out2               => s_out2(4,60),
			lock_lower_row_out => s_locks_lower_out(4,60),
			lock_lower_row_in  => s_locks_lower_in(4,60),
			in1                => s_in1(4,60),
			in2                => (others => '0'),
			lock_row           => s_locks(4),
			piv_found          => s_piv_found,
			row_data           => s_row_data(4),
			col_data           => s_col_data(60)
		);
	s_in1(4,60)            <= s_out1(5,60);
	s_locks_lower_in(4,60) <= s_locks_lower_out(5,60);

		normal_cell_5_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,1),
			fetch              => s_fetch(5,1),
			data_in            => s_data_in(5,1),
			data_out           => s_data_out(5,1),
			out1               => s_out1(5,1),
			out2               => s_out2(5,1),
			lock_lower_row_out => s_locks_lower_out(5,1),
			lock_lower_row_in  => s_locks_lower_in(5,1),
			in1                => s_in1(5,1),
			in2                => s_in2(5,1),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(1)
		);
	s_in1(5,1)            <= s_out1(6,1);
	s_in2(5,1)            <= s_out2(6,2);
	s_locks_lower_in(5,1) <= s_locks_lower_out(6,1);

		normal_cell_5_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,2),
			fetch              => s_fetch(5,2),
			data_in            => s_data_in(5,2),
			data_out           => s_data_out(5,2),
			out1               => s_out1(5,2),
			out2               => s_out2(5,2),
			lock_lower_row_out => s_locks_lower_out(5,2),
			lock_lower_row_in  => s_locks_lower_in(5,2),
			in1                => s_in1(5,2),
			in2                => s_in2(5,2),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(2)
		);
	s_in1(5,2)            <= s_out1(6,2);
	s_in2(5,2)            <= s_out2(6,3);
	s_locks_lower_in(5,2) <= s_locks_lower_out(6,2);

		normal_cell_5_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,3),
			fetch              => s_fetch(5,3),
			data_in            => s_data_in(5,3),
			data_out           => s_data_out(5,3),
			out1               => s_out1(5,3),
			out2               => s_out2(5,3),
			lock_lower_row_out => s_locks_lower_out(5,3),
			lock_lower_row_in  => s_locks_lower_in(5,3),
			in1                => s_in1(5,3),
			in2                => s_in2(5,3),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(3)
		);
	s_in1(5,3)            <= s_out1(6,3);
	s_in2(5,3)            <= s_out2(6,4);
	s_locks_lower_in(5,3) <= s_locks_lower_out(6,3);

		normal_cell_5_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,4),
			fetch              => s_fetch(5,4),
			data_in            => s_data_in(5,4),
			data_out           => s_data_out(5,4),
			out1               => s_out1(5,4),
			out2               => s_out2(5,4),
			lock_lower_row_out => s_locks_lower_out(5,4),
			lock_lower_row_in  => s_locks_lower_in(5,4),
			in1                => s_in1(5,4),
			in2                => s_in2(5,4),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(4)
		);
	s_in1(5,4)            <= s_out1(6,4);
	s_in2(5,4)            <= s_out2(6,5);
	s_locks_lower_in(5,4) <= s_locks_lower_out(6,4);

		normal_cell_5_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,5),
			fetch              => s_fetch(5,5),
			data_in            => s_data_in(5,5),
			data_out           => s_data_out(5,5),
			out1               => s_out1(5,5),
			out2               => s_out2(5,5),
			lock_lower_row_out => s_locks_lower_out(5,5),
			lock_lower_row_in  => s_locks_lower_in(5,5),
			in1                => s_in1(5,5),
			in2                => s_in2(5,5),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(5)
		);
	s_in1(5,5)            <= s_out1(6,5);
	s_in2(5,5)            <= s_out2(6,6);
	s_locks_lower_in(5,5) <= s_locks_lower_out(6,5);

		normal_cell_5_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,6),
			fetch              => s_fetch(5,6),
			data_in            => s_data_in(5,6),
			data_out           => s_data_out(5,6),
			out1               => s_out1(5,6),
			out2               => s_out2(5,6),
			lock_lower_row_out => s_locks_lower_out(5,6),
			lock_lower_row_in  => s_locks_lower_in(5,6),
			in1                => s_in1(5,6),
			in2                => s_in2(5,6),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(6)
		);
	s_in1(5,6)            <= s_out1(6,6);
	s_in2(5,6)            <= s_out2(6,7);
	s_locks_lower_in(5,6) <= s_locks_lower_out(6,6);

		normal_cell_5_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,7),
			fetch              => s_fetch(5,7),
			data_in            => s_data_in(5,7),
			data_out           => s_data_out(5,7),
			out1               => s_out1(5,7),
			out2               => s_out2(5,7),
			lock_lower_row_out => s_locks_lower_out(5,7),
			lock_lower_row_in  => s_locks_lower_in(5,7),
			in1                => s_in1(5,7),
			in2                => s_in2(5,7),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(7)
		);
	s_in1(5,7)            <= s_out1(6,7);
	s_in2(5,7)            <= s_out2(6,8);
	s_locks_lower_in(5,7) <= s_locks_lower_out(6,7);

		normal_cell_5_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,8),
			fetch              => s_fetch(5,8),
			data_in            => s_data_in(5,8),
			data_out           => s_data_out(5,8),
			out1               => s_out1(5,8),
			out2               => s_out2(5,8),
			lock_lower_row_out => s_locks_lower_out(5,8),
			lock_lower_row_in  => s_locks_lower_in(5,8),
			in1                => s_in1(5,8),
			in2                => s_in2(5,8),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(8)
		);
	s_in1(5,8)            <= s_out1(6,8);
	s_in2(5,8)            <= s_out2(6,9);
	s_locks_lower_in(5,8) <= s_locks_lower_out(6,8);

		normal_cell_5_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,9),
			fetch              => s_fetch(5,9),
			data_in            => s_data_in(5,9),
			data_out           => s_data_out(5,9),
			out1               => s_out1(5,9),
			out2               => s_out2(5,9),
			lock_lower_row_out => s_locks_lower_out(5,9),
			lock_lower_row_in  => s_locks_lower_in(5,9),
			in1                => s_in1(5,9),
			in2                => s_in2(5,9),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(9)
		);
	s_in1(5,9)            <= s_out1(6,9);
	s_in2(5,9)            <= s_out2(6,10);
	s_locks_lower_in(5,9) <= s_locks_lower_out(6,9);

		normal_cell_5_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,10),
			fetch              => s_fetch(5,10),
			data_in            => s_data_in(5,10),
			data_out           => s_data_out(5,10),
			out1               => s_out1(5,10),
			out2               => s_out2(5,10),
			lock_lower_row_out => s_locks_lower_out(5,10),
			lock_lower_row_in  => s_locks_lower_in(5,10),
			in1                => s_in1(5,10),
			in2                => s_in2(5,10),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(10)
		);
	s_in1(5,10)            <= s_out1(6,10);
	s_in2(5,10)            <= s_out2(6,11);
	s_locks_lower_in(5,10) <= s_locks_lower_out(6,10);

		normal_cell_5_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,11),
			fetch              => s_fetch(5,11),
			data_in            => s_data_in(5,11),
			data_out           => s_data_out(5,11),
			out1               => s_out1(5,11),
			out2               => s_out2(5,11),
			lock_lower_row_out => s_locks_lower_out(5,11),
			lock_lower_row_in  => s_locks_lower_in(5,11),
			in1                => s_in1(5,11),
			in2                => s_in2(5,11),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(11)
		);
	s_in1(5,11)            <= s_out1(6,11);
	s_in2(5,11)            <= s_out2(6,12);
	s_locks_lower_in(5,11) <= s_locks_lower_out(6,11);

		normal_cell_5_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,12),
			fetch              => s_fetch(5,12),
			data_in            => s_data_in(5,12),
			data_out           => s_data_out(5,12),
			out1               => s_out1(5,12),
			out2               => s_out2(5,12),
			lock_lower_row_out => s_locks_lower_out(5,12),
			lock_lower_row_in  => s_locks_lower_in(5,12),
			in1                => s_in1(5,12),
			in2                => s_in2(5,12),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(12)
		);
	s_in1(5,12)            <= s_out1(6,12);
	s_in2(5,12)            <= s_out2(6,13);
	s_locks_lower_in(5,12) <= s_locks_lower_out(6,12);

		normal_cell_5_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,13),
			fetch              => s_fetch(5,13),
			data_in            => s_data_in(5,13),
			data_out           => s_data_out(5,13),
			out1               => s_out1(5,13),
			out2               => s_out2(5,13),
			lock_lower_row_out => s_locks_lower_out(5,13),
			lock_lower_row_in  => s_locks_lower_in(5,13),
			in1                => s_in1(5,13),
			in2                => s_in2(5,13),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(13)
		);
	s_in1(5,13)            <= s_out1(6,13);
	s_in2(5,13)            <= s_out2(6,14);
	s_locks_lower_in(5,13) <= s_locks_lower_out(6,13);

		normal_cell_5_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,14),
			fetch              => s_fetch(5,14),
			data_in            => s_data_in(5,14),
			data_out           => s_data_out(5,14),
			out1               => s_out1(5,14),
			out2               => s_out2(5,14),
			lock_lower_row_out => s_locks_lower_out(5,14),
			lock_lower_row_in  => s_locks_lower_in(5,14),
			in1                => s_in1(5,14),
			in2                => s_in2(5,14),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(14)
		);
	s_in1(5,14)            <= s_out1(6,14);
	s_in2(5,14)            <= s_out2(6,15);
	s_locks_lower_in(5,14) <= s_locks_lower_out(6,14);

		normal_cell_5_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,15),
			fetch              => s_fetch(5,15),
			data_in            => s_data_in(5,15),
			data_out           => s_data_out(5,15),
			out1               => s_out1(5,15),
			out2               => s_out2(5,15),
			lock_lower_row_out => s_locks_lower_out(5,15),
			lock_lower_row_in  => s_locks_lower_in(5,15),
			in1                => s_in1(5,15),
			in2                => s_in2(5,15),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(15)
		);
	s_in1(5,15)            <= s_out1(6,15);
	s_in2(5,15)            <= s_out2(6,16);
	s_locks_lower_in(5,15) <= s_locks_lower_out(6,15);

		normal_cell_5_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,16),
			fetch              => s_fetch(5,16),
			data_in            => s_data_in(5,16),
			data_out           => s_data_out(5,16),
			out1               => s_out1(5,16),
			out2               => s_out2(5,16),
			lock_lower_row_out => s_locks_lower_out(5,16),
			lock_lower_row_in  => s_locks_lower_in(5,16),
			in1                => s_in1(5,16),
			in2                => s_in2(5,16),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(16)
		);
	s_in1(5,16)            <= s_out1(6,16);
	s_in2(5,16)            <= s_out2(6,17);
	s_locks_lower_in(5,16) <= s_locks_lower_out(6,16);

		normal_cell_5_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,17),
			fetch              => s_fetch(5,17),
			data_in            => s_data_in(5,17),
			data_out           => s_data_out(5,17),
			out1               => s_out1(5,17),
			out2               => s_out2(5,17),
			lock_lower_row_out => s_locks_lower_out(5,17),
			lock_lower_row_in  => s_locks_lower_in(5,17),
			in1                => s_in1(5,17),
			in2                => s_in2(5,17),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(17)
		);
	s_in1(5,17)            <= s_out1(6,17);
	s_in2(5,17)            <= s_out2(6,18);
	s_locks_lower_in(5,17) <= s_locks_lower_out(6,17);

		normal_cell_5_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,18),
			fetch              => s_fetch(5,18),
			data_in            => s_data_in(5,18),
			data_out           => s_data_out(5,18),
			out1               => s_out1(5,18),
			out2               => s_out2(5,18),
			lock_lower_row_out => s_locks_lower_out(5,18),
			lock_lower_row_in  => s_locks_lower_in(5,18),
			in1                => s_in1(5,18),
			in2                => s_in2(5,18),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(18)
		);
	s_in1(5,18)            <= s_out1(6,18);
	s_in2(5,18)            <= s_out2(6,19);
	s_locks_lower_in(5,18) <= s_locks_lower_out(6,18);

		normal_cell_5_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,19),
			fetch              => s_fetch(5,19),
			data_in            => s_data_in(5,19),
			data_out           => s_data_out(5,19),
			out1               => s_out1(5,19),
			out2               => s_out2(5,19),
			lock_lower_row_out => s_locks_lower_out(5,19),
			lock_lower_row_in  => s_locks_lower_in(5,19),
			in1                => s_in1(5,19),
			in2                => s_in2(5,19),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(19)
		);
	s_in1(5,19)            <= s_out1(6,19);
	s_in2(5,19)            <= s_out2(6,20);
	s_locks_lower_in(5,19) <= s_locks_lower_out(6,19);

		normal_cell_5_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,20),
			fetch              => s_fetch(5,20),
			data_in            => s_data_in(5,20),
			data_out           => s_data_out(5,20),
			out1               => s_out1(5,20),
			out2               => s_out2(5,20),
			lock_lower_row_out => s_locks_lower_out(5,20),
			lock_lower_row_in  => s_locks_lower_in(5,20),
			in1                => s_in1(5,20),
			in2                => s_in2(5,20),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(20)
		);
	s_in1(5,20)            <= s_out1(6,20);
	s_in2(5,20)            <= s_out2(6,21);
	s_locks_lower_in(5,20) <= s_locks_lower_out(6,20);

		normal_cell_5_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,21),
			fetch              => s_fetch(5,21),
			data_in            => s_data_in(5,21),
			data_out           => s_data_out(5,21),
			out1               => s_out1(5,21),
			out2               => s_out2(5,21),
			lock_lower_row_out => s_locks_lower_out(5,21),
			lock_lower_row_in  => s_locks_lower_in(5,21),
			in1                => s_in1(5,21),
			in2                => s_in2(5,21),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(21)
		);
	s_in1(5,21)            <= s_out1(6,21);
	s_in2(5,21)            <= s_out2(6,22);
	s_locks_lower_in(5,21) <= s_locks_lower_out(6,21);

		normal_cell_5_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,22),
			fetch              => s_fetch(5,22),
			data_in            => s_data_in(5,22),
			data_out           => s_data_out(5,22),
			out1               => s_out1(5,22),
			out2               => s_out2(5,22),
			lock_lower_row_out => s_locks_lower_out(5,22),
			lock_lower_row_in  => s_locks_lower_in(5,22),
			in1                => s_in1(5,22),
			in2                => s_in2(5,22),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(22)
		);
	s_in1(5,22)            <= s_out1(6,22);
	s_in2(5,22)            <= s_out2(6,23);
	s_locks_lower_in(5,22) <= s_locks_lower_out(6,22);

		normal_cell_5_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,23),
			fetch              => s_fetch(5,23),
			data_in            => s_data_in(5,23),
			data_out           => s_data_out(5,23),
			out1               => s_out1(5,23),
			out2               => s_out2(5,23),
			lock_lower_row_out => s_locks_lower_out(5,23),
			lock_lower_row_in  => s_locks_lower_in(5,23),
			in1                => s_in1(5,23),
			in2                => s_in2(5,23),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(23)
		);
	s_in1(5,23)            <= s_out1(6,23);
	s_in2(5,23)            <= s_out2(6,24);
	s_locks_lower_in(5,23) <= s_locks_lower_out(6,23);

		normal_cell_5_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,24),
			fetch              => s_fetch(5,24),
			data_in            => s_data_in(5,24),
			data_out           => s_data_out(5,24),
			out1               => s_out1(5,24),
			out2               => s_out2(5,24),
			lock_lower_row_out => s_locks_lower_out(5,24),
			lock_lower_row_in  => s_locks_lower_in(5,24),
			in1                => s_in1(5,24),
			in2                => s_in2(5,24),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(24)
		);
	s_in1(5,24)            <= s_out1(6,24);
	s_in2(5,24)            <= s_out2(6,25);
	s_locks_lower_in(5,24) <= s_locks_lower_out(6,24);

		normal_cell_5_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,25),
			fetch              => s_fetch(5,25),
			data_in            => s_data_in(5,25),
			data_out           => s_data_out(5,25),
			out1               => s_out1(5,25),
			out2               => s_out2(5,25),
			lock_lower_row_out => s_locks_lower_out(5,25),
			lock_lower_row_in  => s_locks_lower_in(5,25),
			in1                => s_in1(5,25),
			in2                => s_in2(5,25),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(25)
		);
	s_in1(5,25)            <= s_out1(6,25);
	s_in2(5,25)            <= s_out2(6,26);
	s_locks_lower_in(5,25) <= s_locks_lower_out(6,25);

		normal_cell_5_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,26),
			fetch              => s_fetch(5,26),
			data_in            => s_data_in(5,26),
			data_out           => s_data_out(5,26),
			out1               => s_out1(5,26),
			out2               => s_out2(5,26),
			lock_lower_row_out => s_locks_lower_out(5,26),
			lock_lower_row_in  => s_locks_lower_in(5,26),
			in1                => s_in1(5,26),
			in2                => s_in2(5,26),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(26)
		);
	s_in1(5,26)            <= s_out1(6,26);
	s_in2(5,26)            <= s_out2(6,27);
	s_locks_lower_in(5,26) <= s_locks_lower_out(6,26);

		normal_cell_5_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,27),
			fetch              => s_fetch(5,27),
			data_in            => s_data_in(5,27),
			data_out           => s_data_out(5,27),
			out1               => s_out1(5,27),
			out2               => s_out2(5,27),
			lock_lower_row_out => s_locks_lower_out(5,27),
			lock_lower_row_in  => s_locks_lower_in(5,27),
			in1                => s_in1(5,27),
			in2                => s_in2(5,27),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(27)
		);
	s_in1(5,27)            <= s_out1(6,27);
	s_in2(5,27)            <= s_out2(6,28);
	s_locks_lower_in(5,27) <= s_locks_lower_out(6,27);

		normal_cell_5_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,28),
			fetch              => s_fetch(5,28),
			data_in            => s_data_in(5,28),
			data_out           => s_data_out(5,28),
			out1               => s_out1(5,28),
			out2               => s_out2(5,28),
			lock_lower_row_out => s_locks_lower_out(5,28),
			lock_lower_row_in  => s_locks_lower_in(5,28),
			in1                => s_in1(5,28),
			in2                => s_in2(5,28),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(28)
		);
	s_in1(5,28)            <= s_out1(6,28);
	s_in2(5,28)            <= s_out2(6,29);
	s_locks_lower_in(5,28) <= s_locks_lower_out(6,28);

		normal_cell_5_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,29),
			fetch              => s_fetch(5,29),
			data_in            => s_data_in(5,29),
			data_out           => s_data_out(5,29),
			out1               => s_out1(5,29),
			out2               => s_out2(5,29),
			lock_lower_row_out => s_locks_lower_out(5,29),
			lock_lower_row_in  => s_locks_lower_in(5,29),
			in1                => s_in1(5,29),
			in2                => s_in2(5,29),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(29)
		);
	s_in1(5,29)            <= s_out1(6,29);
	s_in2(5,29)            <= s_out2(6,30);
	s_locks_lower_in(5,29) <= s_locks_lower_out(6,29);

		normal_cell_5_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,30),
			fetch              => s_fetch(5,30),
			data_in            => s_data_in(5,30),
			data_out           => s_data_out(5,30),
			out1               => s_out1(5,30),
			out2               => s_out2(5,30),
			lock_lower_row_out => s_locks_lower_out(5,30),
			lock_lower_row_in  => s_locks_lower_in(5,30),
			in1                => s_in1(5,30),
			in2                => s_in2(5,30),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(30)
		);
	s_in1(5,30)            <= s_out1(6,30);
	s_in2(5,30)            <= s_out2(6,31);
	s_locks_lower_in(5,30) <= s_locks_lower_out(6,30);

		normal_cell_5_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,31),
			fetch              => s_fetch(5,31),
			data_in            => s_data_in(5,31),
			data_out           => s_data_out(5,31),
			out1               => s_out1(5,31),
			out2               => s_out2(5,31),
			lock_lower_row_out => s_locks_lower_out(5,31),
			lock_lower_row_in  => s_locks_lower_in(5,31),
			in1                => s_in1(5,31),
			in2                => s_in2(5,31),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(31)
		);
	s_in1(5,31)            <= s_out1(6,31);
	s_in2(5,31)            <= s_out2(6,32);
	s_locks_lower_in(5,31) <= s_locks_lower_out(6,31);

		normal_cell_5_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,32),
			fetch              => s_fetch(5,32),
			data_in            => s_data_in(5,32),
			data_out           => s_data_out(5,32),
			out1               => s_out1(5,32),
			out2               => s_out2(5,32),
			lock_lower_row_out => s_locks_lower_out(5,32),
			lock_lower_row_in  => s_locks_lower_in(5,32),
			in1                => s_in1(5,32),
			in2                => s_in2(5,32),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(32)
		);
	s_in1(5,32)            <= s_out1(6,32);
	s_in2(5,32)            <= s_out2(6,33);
	s_locks_lower_in(5,32) <= s_locks_lower_out(6,32);

		normal_cell_5_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,33),
			fetch              => s_fetch(5,33),
			data_in            => s_data_in(5,33),
			data_out           => s_data_out(5,33),
			out1               => s_out1(5,33),
			out2               => s_out2(5,33),
			lock_lower_row_out => s_locks_lower_out(5,33),
			lock_lower_row_in  => s_locks_lower_in(5,33),
			in1                => s_in1(5,33),
			in2                => s_in2(5,33),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(33)
		);
	s_in1(5,33)            <= s_out1(6,33);
	s_in2(5,33)            <= s_out2(6,34);
	s_locks_lower_in(5,33) <= s_locks_lower_out(6,33);

		normal_cell_5_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,34),
			fetch              => s_fetch(5,34),
			data_in            => s_data_in(5,34),
			data_out           => s_data_out(5,34),
			out1               => s_out1(5,34),
			out2               => s_out2(5,34),
			lock_lower_row_out => s_locks_lower_out(5,34),
			lock_lower_row_in  => s_locks_lower_in(5,34),
			in1                => s_in1(5,34),
			in2                => s_in2(5,34),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(34)
		);
	s_in1(5,34)            <= s_out1(6,34);
	s_in2(5,34)            <= s_out2(6,35);
	s_locks_lower_in(5,34) <= s_locks_lower_out(6,34);

		normal_cell_5_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,35),
			fetch              => s_fetch(5,35),
			data_in            => s_data_in(5,35),
			data_out           => s_data_out(5,35),
			out1               => s_out1(5,35),
			out2               => s_out2(5,35),
			lock_lower_row_out => s_locks_lower_out(5,35),
			lock_lower_row_in  => s_locks_lower_in(5,35),
			in1                => s_in1(5,35),
			in2                => s_in2(5,35),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(35)
		);
	s_in1(5,35)            <= s_out1(6,35);
	s_in2(5,35)            <= s_out2(6,36);
	s_locks_lower_in(5,35) <= s_locks_lower_out(6,35);

		normal_cell_5_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,36),
			fetch              => s_fetch(5,36),
			data_in            => s_data_in(5,36),
			data_out           => s_data_out(5,36),
			out1               => s_out1(5,36),
			out2               => s_out2(5,36),
			lock_lower_row_out => s_locks_lower_out(5,36),
			lock_lower_row_in  => s_locks_lower_in(5,36),
			in1                => s_in1(5,36),
			in2                => s_in2(5,36),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(36)
		);
	s_in1(5,36)            <= s_out1(6,36);
	s_in2(5,36)            <= s_out2(6,37);
	s_locks_lower_in(5,36) <= s_locks_lower_out(6,36);

		normal_cell_5_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,37),
			fetch              => s_fetch(5,37),
			data_in            => s_data_in(5,37),
			data_out           => s_data_out(5,37),
			out1               => s_out1(5,37),
			out2               => s_out2(5,37),
			lock_lower_row_out => s_locks_lower_out(5,37),
			lock_lower_row_in  => s_locks_lower_in(5,37),
			in1                => s_in1(5,37),
			in2                => s_in2(5,37),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(37)
		);
	s_in1(5,37)            <= s_out1(6,37);
	s_in2(5,37)            <= s_out2(6,38);
	s_locks_lower_in(5,37) <= s_locks_lower_out(6,37);

		normal_cell_5_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,38),
			fetch              => s_fetch(5,38),
			data_in            => s_data_in(5,38),
			data_out           => s_data_out(5,38),
			out1               => s_out1(5,38),
			out2               => s_out2(5,38),
			lock_lower_row_out => s_locks_lower_out(5,38),
			lock_lower_row_in  => s_locks_lower_in(5,38),
			in1                => s_in1(5,38),
			in2                => s_in2(5,38),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(38)
		);
	s_in1(5,38)            <= s_out1(6,38);
	s_in2(5,38)            <= s_out2(6,39);
	s_locks_lower_in(5,38) <= s_locks_lower_out(6,38);

		normal_cell_5_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,39),
			fetch              => s_fetch(5,39),
			data_in            => s_data_in(5,39),
			data_out           => s_data_out(5,39),
			out1               => s_out1(5,39),
			out2               => s_out2(5,39),
			lock_lower_row_out => s_locks_lower_out(5,39),
			lock_lower_row_in  => s_locks_lower_in(5,39),
			in1                => s_in1(5,39),
			in2                => s_in2(5,39),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(39)
		);
	s_in1(5,39)            <= s_out1(6,39);
	s_in2(5,39)            <= s_out2(6,40);
	s_locks_lower_in(5,39) <= s_locks_lower_out(6,39);

		normal_cell_5_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,40),
			fetch              => s_fetch(5,40),
			data_in            => s_data_in(5,40),
			data_out           => s_data_out(5,40),
			out1               => s_out1(5,40),
			out2               => s_out2(5,40),
			lock_lower_row_out => s_locks_lower_out(5,40),
			lock_lower_row_in  => s_locks_lower_in(5,40),
			in1                => s_in1(5,40),
			in2                => s_in2(5,40),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(40)
		);
	s_in1(5,40)            <= s_out1(6,40);
	s_in2(5,40)            <= s_out2(6,41);
	s_locks_lower_in(5,40) <= s_locks_lower_out(6,40);

		normal_cell_5_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,41),
			fetch              => s_fetch(5,41),
			data_in            => s_data_in(5,41),
			data_out           => s_data_out(5,41),
			out1               => s_out1(5,41),
			out2               => s_out2(5,41),
			lock_lower_row_out => s_locks_lower_out(5,41),
			lock_lower_row_in  => s_locks_lower_in(5,41),
			in1                => s_in1(5,41),
			in2                => s_in2(5,41),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(41)
		);
	s_in1(5,41)            <= s_out1(6,41);
	s_in2(5,41)            <= s_out2(6,42);
	s_locks_lower_in(5,41) <= s_locks_lower_out(6,41);

		normal_cell_5_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,42),
			fetch              => s_fetch(5,42),
			data_in            => s_data_in(5,42),
			data_out           => s_data_out(5,42),
			out1               => s_out1(5,42),
			out2               => s_out2(5,42),
			lock_lower_row_out => s_locks_lower_out(5,42),
			lock_lower_row_in  => s_locks_lower_in(5,42),
			in1                => s_in1(5,42),
			in2                => s_in2(5,42),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(42)
		);
	s_in1(5,42)            <= s_out1(6,42);
	s_in2(5,42)            <= s_out2(6,43);
	s_locks_lower_in(5,42) <= s_locks_lower_out(6,42);

		normal_cell_5_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,43),
			fetch              => s_fetch(5,43),
			data_in            => s_data_in(5,43),
			data_out           => s_data_out(5,43),
			out1               => s_out1(5,43),
			out2               => s_out2(5,43),
			lock_lower_row_out => s_locks_lower_out(5,43),
			lock_lower_row_in  => s_locks_lower_in(5,43),
			in1                => s_in1(5,43),
			in2                => s_in2(5,43),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(43)
		);
	s_in1(5,43)            <= s_out1(6,43);
	s_in2(5,43)            <= s_out2(6,44);
	s_locks_lower_in(5,43) <= s_locks_lower_out(6,43);

		normal_cell_5_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,44),
			fetch              => s_fetch(5,44),
			data_in            => s_data_in(5,44),
			data_out           => s_data_out(5,44),
			out1               => s_out1(5,44),
			out2               => s_out2(5,44),
			lock_lower_row_out => s_locks_lower_out(5,44),
			lock_lower_row_in  => s_locks_lower_in(5,44),
			in1                => s_in1(5,44),
			in2                => s_in2(5,44),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(44)
		);
	s_in1(5,44)            <= s_out1(6,44);
	s_in2(5,44)            <= s_out2(6,45);
	s_locks_lower_in(5,44) <= s_locks_lower_out(6,44);

		normal_cell_5_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,45),
			fetch              => s_fetch(5,45),
			data_in            => s_data_in(5,45),
			data_out           => s_data_out(5,45),
			out1               => s_out1(5,45),
			out2               => s_out2(5,45),
			lock_lower_row_out => s_locks_lower_out(5,45),
			lock_lower_row_in  => s_locks_lower_in(5,45),
			in1                => s_in1(5,45),
			in2                => s_in2(5,45),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(45)
		);
	s_in1(5,45)            <= s_out1(6,45);
	s_in2(5,45)            <= s_out2(6,46);
	s_locks_lower_in(5,45) <= s_locks_lower_out(6,45);

		normal_cell_5_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,46),
			fetch              => s_fetch(5,46),
			data_in            => s_data_in(5,46),
			data_out           => s_data_out(5,46),
			out1               => s_out1(5,46),
			out2               => s_out2(5,46),
			lock_lower_row_out => s_locks_lower_out(5,46),
			lock_lower_row_in  => s_locks_lower_in(5,46),
			in1                => s_in1(5,46),
			in2                => s_in2(5,46),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(46)
		);
	s_in1(5,46)            <= s_out1(6,46);
	s_in2(5,46)            <= s_out2(6,47);
	s_locks_lower_in(5,46) <= s_locks_lower_out(6,46);

		normal_cell_5_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,47),
			fetch              => s_fetch(5,47),
			data_in            => s_data_in(5,47),
			data_out           => s_data_out(5,47),
			out1               => s_out1(5,47),
			out2               => s_out2(5,47),
			lock_lower_row_out => s_locks_lower_out(5,47),
			lock_lower_row_in  => s_locks_lower_in(5,47),
			in1                => s_in1(5,47),
			in2                => s_in2(5,47),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(47)
		);
	s_in1(5,47)            <= s_out1(6,47);
	s_in2(5,47)            <= s_out2(6,48);
	s_locks_lower_in(5,47) <= s_locks_lower_out(6,47);

		normal_cell_5_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,48),
			fetch              => s_fetch(5,48),
			data_in            => s_data_in(5,48),
			data_out           => s_data_out(5,48),
			out1               => s_out1(5,48),
			out2               => s_out2(5,48),
			lock_lower_row_out => s_locks_lower_out(5,48),
			lock_lower_row_in  => s_locks_lower_in(5,48),
			in1                => s_in1(5,48),
			in2                => s_in2(5,48),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(48)
		);
	s_in1(5,48)            <= s_out1(6,48);
	s_in2(5,48)            <= s_out2(6,49);
	s_locks_lower_in(5,48) <= s_locks_lower_out(6,48);

		normal_cell_5_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,49),
			fetch              => s_fetch(5,49),
			data_in            => s_data_in(5,49),
			data_out           => s_data_out(5,49),
			out1               => s_out1(5,49),
			out2               => s_out2(5,49),
			lock_lower_row_out => s_locks_lower_out(5,49),
			lock_lower_row_in  => s_locks_lower_in(5,49),
			in1                => s_in1(5,49),
			in2                => s_in2(5,49),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(49)
		);
	s_in1(5,49)            <= s_out1(6,49);
	s_in2(5,49)            <= s_out2(6,50);
	s_locks_lower_in(5,49) <= s_locks_lower_out(6,49);

		normal_cell_5_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,50),
			fetch              => s_fetch(5,50),
			data_in            => s_data_in(5,50),
			data_out           => s_data_out(5,50),
			out1               => s_out1(5,50),
			out2               => s_out2(5,50),
			lock_lower_row_out => s_locks_lower_out(5,50),
			lock_lower_row_in  => s_locks_lower_in(5,50),
			in1                => s_in1(5,50),
			in2                => s_in2(5,50),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(50)
		);
	s_in1(5,50)            <= s_out1(6,50);
	s_in2(5,50)            <= s_out2(6,51);
	s_locks_lower_in(5,50) <= s_locks_lower_out(6,50);

		normal_cell_5_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,51),
			fetch              => s_fetch(5,51),
			data_in            => s_data_in(5,51),
			data_out           => s_data_out(5,51),
			out1               => s_out1(5,51),
			out2               => s_out2(5,51),
			lock_lower_row_out => s_locks_lower_out(5,51),
			lock_lower_row_in  => s_locks_lower_in(5,51),
			in1                => s_in1(5,51),
			in2                => s_in2(5,51),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(51)
		);
	s_in1(5,51)            <= s_out1(6,51);
	s_in2(5,51)            <= s_out2(6,52);
	s_locks_lower_in(5,51) <= s_locks_lower_out(6,51);

		normal_cell_5_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,52),
			fetch              => s_fetch(5,52),
			data_in            => s_data_in(5,52),
			data_out           => s_data_out(5,52),
			out1               => s_out1(5,52),
			out2               => s_out2(5,52),
			lock_lower_row_out => s_locks_lower_out(5,52),
			lock_lower_row_in  => s_locks_lower_in(5,52),
			in1                => s_in1(5,52),
			in2                => s_in2(5,52),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(52)
		);
	s_in1(5,52)            <= s_out1(6,52);
	s_in2(5,52)            <= s_out2(6,53);
	s_locks_lower_in(5,52) <= s_locks_lower_out(6,52);

		normal_cell_5_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,53),
			fetch              => s_fetch(5,53),
			data_in            => s_data_in(5,53),
			data_out           => s_data_out(5,53),
			out1               => s_out1(5,53),
			out2               => s_out2(5,53),
			lock_lower_row_out => s_locks_lower_out(5,53),
			lock_lower_row_in  => s_locks_lower_in(5,53),
			in1                => s_in1(5,53),
			in2                => s_in2(5,53),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(53)
		);
	s_in1(5,53)            <= s_out1(6,53);
	s_in2(5,53)            <= s_out2(6,54);
	s_locks_lower_in(5,53) <= s_locks_lower_out(6,53);

		normal_cell_5_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,54),
			fetch              => s_fetch(5,54),
			data_in            => s_data_in(5,54),
			data_out           => s_data_out(5,54),
			out1               => s_out1(5,54),
			out2               => s_out2(5,54),
			lock_lower_row_out => s_locks_lower_out(5,54),
			lock_lower_row_in  => s_locks_lower_in(5,54),
			in1                => s_in1(5,54),
			in2                => s_in2(5,54),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(54)
		);
	s_in1(5,54)            <= s_out1(6,54);
	s_in2(5,54)            <= s_out2(6,55);
	s_locks_lower_in(5,54) <= s_locks_lower_out(6,54);

		normal_cell_5_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,55),
			fetch              => s_fetch(5,55),
			data_in            => s_data_in(5,55),
			data_out           => s_data_out(5,55),
			out1               => s_out1(5,55),
			out2               => s_out2(5,55),
			lock_lower_row_out => s_locks_lower_out(5,55),
			lock_lower_row_in  => s_locks_lower_in(5,55),
			in1                => s_in1(5,55),
			in2                => s_in2(5,55),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(55)
		);
	s_in1(5,55)            <= s_out1(6,55);
	s_in2(5,55)            <= s_out2(6,56);
	s_locks_lower_in(5,55) <= s_locks_lower_out(6,55);

		normal_cell_5_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,56),
			fetch              => s_fetch(5,56),
			data_in            => s_data_in(5,56),
			data_out           => s_data_out(5,56),
			out1               => s_out1(5,56),
			out2               => s_out2(5,56),
			lock_lower_row_out => s_locks_lower_out(5,56),
			lock_lower_row_in  => s_locks_lower_in(5,56),
			in1                => s_in1(5,56),
			in2                => s_in2(5,56),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(56)
		);
	s_in1(5,56)            <= s_out1(6,56);
	s_in2(5,56)            <= s_out2(6,57);
	s_locks_lower_in(5,56) <= s_locks_lower_out(6,56);

		normal_cell_5_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,57),
			fetch              => s_fetch(5,57),
			data_in            => s_data_in(5,57),
			data_out           => s_data_out(5,57),
			out1               => s_out1(5,57),
			out2               => s_out2(5,57),
			lock_lower_row_out => s_locks_lower_out(5,57),
			lock_lower_row_in  => s_locks_lower_in(5,57),
			in1                => s_in1(5,57),
			in2                => s_in2(5,57),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(57)
		);
	s_in1(5,57)            <= s_out1(6,57);
	s_in2(5,57)            <= s_out2(6,58);
	s_locks_lower_in(5,57) <= s_locks_lower_out(6,57);

		normal_cell_5_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,58),
			fetch              => s_fetch(5,58),
			data_in            => s_data_in(5,58),
			data_out           => s_data_out(5,58),
			out1               => s_out1(5,58),
			out2               => s_out2(5,58),
			lock_lower_row_out => s_locks_lower_out(5,58),
			lock_lower_row_in  => s_locks_lower_in(5,58),
			in1                => s_in1(5,58),
			in2                => s_in2(5,58),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(58)
		);
	s_in1(5,58)            <= s_out1(6,58);
	s_in2(5,58)            <= s_out2(6,59);
	s_locks_lower_in(5,58) <= s_locks_lower_out(6,58);

		normal_cell_5_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,59),
			fetch              => s_fetch(5,59),
			data_in            => s_data_in(5,59),
			data_out           => s_data_out(5,59),
			out1               => s_out1(5,59),
			out2               => s_out2(5,59),
			lock_lower_row_out => s_locks_lower_out(5,59),
			lock_lower_row_in  => s_locks_lower_in(5,59),
			in1                => s_in1(5,59),
			in2                => s_in2(5,59),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(59)
		);
	s_in1(5,59)            <= s_out1(6,59);
	s_in2(5,59)            <= s_out2(6,60);
	s_locks_lower_in(5,59) <= s_locks_lower_out(6,59);

		last_col_cell_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(5,60),
			fetch              => s_fetch(5,60),
			data_in            => s_data_in(5,60),
			data_out           => s_data_out(5,60),
			out1               => s_out1(5,60),
			out2               => s_out2(5,60),
			lock_lower_row_out => s_locks_lower_out(5,60),
			lock_lower_row_in  => s_locks_lower_in(5,60),
			in1                => s_in1(5,60),
			in2                => (others => '0'),
			lock_row           => s_locks(5),
			piv_found          => s_piv_found,
			row_data           => s_row_data(5),
			col_data           => s_col_data(60)
		);
	s_in1(5,60)            <= s_out1(6,60);
	s_locks_lower_in(5,60) <= s_locks_lower_out(6,60);

		normal_cell_6_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,1),
			fetch              => s_fetch(6,1),
			data_in            => s_data_in(6,1),
			data_out           => s_data_out(6,1),
			out1               => s_out1(6,1),
			out2               => s_out2(6,1),
			lock_lower_row_out => s_locks_lower_out(6,1),
			lock_lower_row_in  => s_locks_lower_in(6,1),
			in1                => s_in1(6,1),
			in2                => s_in2(6,1),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(1)
		);
	s_in1(6,1)            <= s_out1(7,1);
	s_in2(6,1)            <= s_out2(7,2);
	s_locks_lower_in(6,1) <= s_locks_lower_out(7,1);

		normal_cell_6_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,2),
			fetch              => s_fetch(6,2),
			data_in            => s_data_in(6,2),
			data_out           => s_data_out(6,2),
			out1               => s_out1(6,2),
			out2               => s_out2(6,2),
			lock_lower_row_out => s_locks_lower_out(6,2),
			lock_lower_row_in  => s_locks_lower_in(6,2),
			in1                => s_in1(6,2),
			in2                => s_in2(6,2),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(2)
		);
	s_in1(6,2)            <= s_out1(7,2);
	s_in2(6,2)            <= s_out2(7,3);
	s_locks_lower_in(6,2) <= s_locks_lower_out(7,2);

		normal_cell_6_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,3),
			fetch              => s_fetch(6,3),
			data_in            => s_data_in(6,3),
			data_out           => s_data_out(6,3),
			out1               => s_out1(6,3),
			out2               => s_out2(6,3),
			lock_lower_row_out => s_locks_lower_out(6,3),
			lock_lower_row_in  => s_locks_lower_in(6,3),
			in1                => s_in1(6,3),
			in2                => s_in2(6,3),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(3)
		);
	s_in1(6,3)            <= s_out1(7,3);
	s_in2(6,3)            <= s_out2(7,4);
	s_locks_lower_in(6,3) <= s_locks_lower_out(7,3);

		normal_cell_6_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,4),
			fetch              => s_fetch(6,4),
			data_in            => s_data_in(6,4),
			data_out           => s_data_out(6,4),
			out1               => s_out1(6,4),
			out2               => s_out2(6,4),
			lock_lower_row_out => s_locks_lower_out(6,4),
			lock_lower_row_in  => s_locks_lower_in(6,4),
			in1                => s_in1(6,4),
			in2                => s_in2(6,4),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(4)
		);
	s_in1(6,4)            <= s_out1(7,4);
	s_in2(6,4)            <= s_out2(7,5);
	s_locks_lower_in(6,4) <= s_locks_lower_out(7,4);

		normal_cell_6_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,5),
			fetch              => s_fetch(6,5),
			data_in            => s_data_in(6,5),
			data_out           => s_data_out(6,5),
			out1               => s_out1(6,5),
			out2               => s_out2(6,5),
			lock_lower_row_out => s_locks_lower_out(6,5),
			lock_lower_row_in  => s_locks_lower_in(6,5),
			in1                => s_in1(6,5),
			in2                => s_in2(6,5),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(5)
		);
	s_in1(6,5)            <= s_out1(7,5);
	s_in2(6,5)            <= s_out2(7,6);
	s_locks_lower_in(6,5) <= s_locks_lower_out(7,5);

		normal_cell_6_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,6),
			fetch              => s_fetch(6,6),
			data_in            => s_data_in(6,6),
			data_out           => s_data_out(6,6),
			out1               => s_out1(6,6),
			out2               => s_out2(6,6),
			lock_lower_row_out => s_locks_lower_out(6,6),
			lock_lower_row_in  => s_locks_lower_in(6,6),
			in1                => s_in1(6,6),
			in2                => s_in2(6,6),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(6)
		);
	s_in1(6,6)            <= s_out1(7,6);
	s_in2(6,6)            <= s_out2(7,7);
	s_locks_lower_in(6,6) <= s_locks_lower_out(7,6);

		normal_cell_6_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,7),
			fetch              => s_fetch(6,7),
			data_in            => s_data_in(6,7),
			data_out           => s_data_out(6,7),
			out1               => s_out1(6,7),
			out2               => s_out2(6,7),
			lock_lower_row_out => s_locks_lower_out(6,7),
			lock_lower_row_in  => s_locks_lower_in(6,7),
			in1                => s_in1(6,7),
			in2                => s_in2(6,7),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(7)
		);
	s_in1(6,7)            <= s_out1(7,7);
	s_in2(6,7)            <= s_out2(7,8);
	s_locks_lower_in(6,7) <= s_locks_lower_out(7,7);

		normal_cell_6_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,8),
			fetch              => s_fetch(6,8),
			data_in            => s_data_in(6,8),
			data_out           => s_data_out(6,8),
			out1               => s_out1(6,8),
			out2               => s_out2(6,8),
			lock_lower_row_out => s_locks_lower_out(6,8),
			lock_lower_row_in  => s_locks_lower_in(6,8),
			in1                => s_in1(6,8),
			in2                => s_in2(6,8),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(8)
		);
	s_in1(6,8)            <= s_out1(7,8);
	s_in2(6,8)            <= s_out2(7,9);
	s_locks_lower_in(6,8) <= s_locks_lower_out(7,8);

		normal_cell_6_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,9),
			fetch              => s_fetch(6,9),
			data_in            => s_data_in(6,9),
			data_out           => s_data_out(6,9),
			out1               => s_out1(6,9),
			out2               => s_out2(6,9),
			lock_lower_row_out => s_locks_lower_out(6,9),
			lock_lower_row_in  => s_locks_lower_in(6,9),
			in1                => s_in1(6,9),
			in2                => s_in2(6,9),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(9)
		);
	s_in1(6,9)            <= s_out1(7,9);
	s_in2(6,9)            <= s_out2(7,10);
	s_locks_lower_in(6,9) <= s_locks_lower_out(7,9);

		normal_cell_6_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,10),
			fetch              => s_fetch(6,10),
			data_in            => s_data_in(6,10),
			data_out           => s_data_out(6,10),
			out1               => s_out1(6,10),
			out2               => s_out2(6,10),
			lock_lower_row_out => s_locks_lower_out(6,10),
			lock_lower_row_in  => s_locks_lower_in(6,10),
			in1                => s_in1(6,10),
			in2                => s_in2(6,10),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(10)
		);
	s_in1(6,10)            <= s_out1(7,10);
	s_in2(6,10)            <= s_out2(7,11);
	s_locks_lower_in(6,10) <= s_locks_lower_out(7,10);

		normal_cell_6_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,11),
			fetch              => s_fetch(6,11),
			data_in            => s_data_in(6,11),
			data_out           => s_data_out(6,11),
			out1               => s_out1(6,11),
			out2               => s_out2(6,11),
			lock_lower_row_out => s_locks_lower_out(6,11),
			lock_lower_row_in  => s_locks_lower_in(6,11),
			in1                => s_in1(6,11),
			in2                => s_in2(6,11),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(11)
		);
	s_in1(6,11)            <= s_out1(7,11);
	s_in2(6,11)            <= s_out2(7,12);
	s_locks_lower_in(6,11) <= s_locks_lower_out(7,11);

		normal_cell_6_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,12),
			fetch              => s_fetch(6,12),
			data_in            => s_data_in(6,12),
			data_out           => s_data_out(6,12),
			out1               => s_out1(6,12),
			out2               => s_out2(6,12),
			lock_lower_row_out => s_locks_lower_out(6,12),
			lock_lower_row_in  => s_locks_lower_in(6,12),
			in1                => s_in1(6,12),
			in2                => s_in2(6,12),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(12)
		);
	s_in1(6,12)            <= s_out1(7,12);
	s_in2(6,12)            <= s_out2(7,13);
	s_locks_lower_in(6,12) <= s_locks_lower_out(7,12);

		normal_cell_6_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,13),
			fetch              => s_fetch(6,13),
			data_in            => s_data_in(6,13),
			data_out           => s_data_out(6,13),
			out1               => s_out1(6,13),
			out2               => s_out2(6,13),
			lock_lower_row_out => s_locks_lower_out(6,13),
			lock_lower_row_in  => s_locks_lower_in(6,13),
			in1                => s_in1(6,13),
			in2                => s_in2(6,13),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(13)
		);
	s_in1(6,13)            <= s_out1(7,13);
	s_in2(6,13)            <= s_out2(7,14);
	s_locks_lower_in(6,13) <= s_locks_lower_out(7,13);

		normal_cell_6_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,14),
			fetch              => s_fetch(6,14),
			data_in            => s_data_in(6,14),
			data_out           => s_data_out(6,14),
			out1               => s_out1(6,14),
			out2               => s_out2(6,14),
			lock_lower_row_out => s_locks_lower_out(6,14),
			lock_lower_row_in  => s_locks_lower_in(6,14),
			in1                => s_in1(6,14),
			in2                => s_in2(6,14),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(14)
		);
	s_in1(6,14)            <= s_out1(7,14);
	s_in2(6,14)            <= s_out2(7,15);
	s_locks_lower_in(6,14) <= s_locks_lower_out(7,14);

		normal_cell_6_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,15),
			fetch              => s_fetch(6,15),
			data_in            => s_data_in(6,15),
			data_out           => s_data_out(6,15),
			out1               => s_out1(6,15),
			out2               => s_out2(6,15),
			lock_lower_row_out => s_locks_lower_out(6,15),
			lock_lower_row_in  => s_locks_lower_in(6,15),
			in1                => s_in1(6,15),
			in2                => s_in2(6,15),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(15)
		);
	s_in1(6,15)            <= s_out1(7,15);
	s_in2(6,15)            <= s_out2(7,16);
	s_locks_lower_in(6,15) <= s_locks_lower_out(7,15);

		normal_cell_6_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,16),
			fetch              => s_fetch(6,16),
			data_in            => s_data_in(6,16),
			data_out           => s_data_out(6,16),
			out1               => s_out1(6,16),
			out2               => s_out2(6,16),
			lock_lower_row_out => s_locks_lower_out(6,16),
			lock_lower_row_in  => s_locks_lower_in(6,16),
			in1                => s_in1(6,16),
			in2                => s_in2(6,16),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(16)
		);
	s_in1(6,16)            <= s_out1(7,16);
	s_in2(6,16)            <= s_out2(7,17);
	s_locks_lower_in(6,16) <= s_locks_lower_out(7,16);

		normal_cell_6_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,17),
			fetch              => s_fetch(6,17),
			data_in            => s_data_in(6,17),
			data_out           => s_data_out(6,17),
			out1               => s_out1(6,17),
			out2               => s_out2(6,17),
			lock_lower_row_out => s_locks_lower_out(6,17),
			lock_lower_row_in  => s_locks_lower_in(6,17),
			in1                => s_in1(6,17),
			in2                => s_in2(6,17),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(17)
		);
	s_in1(6,17)            <= s_out1(7,17);
	s_in2(6,17)            <= s_out2(7,18);
	s_locks_lower_in(6,17) <= s_locks_lower_out(7,17);

		normal_cell_6_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,18),
			fetch              => s_fetch(6,18),
			data_in            => s_data_in(6,18),
			data_out           => s_data_out(6,18),
			out1               => s_out1(6,18),
			out2               => s_out2(6,18),
			lock_lower_row_out => s_locks_lower_out(6,18),
			lock_lower_row_in  => s_locks_lower_in(6,18),
			in1                => s_in1(6,18),
			in2                => s_in2(6,18),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(18)
		);
	s_in1(6,18)            <= s_out1(7,18);
	s_in2(6,18)            <= s_out2(7,19);
	s_locks_lower_in(6,18) <= s_locks_lower_out(7,18);

		normal_cell_6_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,19),
			fetch              => s_fetch(6,19),
			data_in            => s_data_in(6,19),
			data_out           => s_data_out(6,19),
			out1               => s_out1(6,19),
			out2               => s_out2(6,19),
			lock_lower_row_out => s_locks_lower_out(6,19),
			lock_lower_row_in  => s_locks_lower_in(6,19),
			in1                => s_in1(6,19),
			in2                => s_in2(6,19),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(19)
		);
	s_in1(6,19)            <= s_out1(7,19);
	s_in2(6,19)            <= s_out2(7,20);
	s_locks_lower_in(6,19) <= s_locks_lower_out(7,19);

		normal_cell_6_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,20),
			fetch              => s_fetch(6,20),
			data_in            => s_data_in(6,20),
			data_out           => s_data_out(6,20),
			out1               => s_out1(6,20),
			out2               => s_out2(6,20),
			lock_lower_row_out => s_locks_lower_out(6,20),
			lock_lower_row_in  => s_locks_lower_in(6,20),
			in1                => s_in1(6,20),
			in2                => s_in2(6,20),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(20)
		);
	s_in1(6,20)            <= s_out1(7,20);
	s_in2(6,20)            <= s_out2(7,21);
	s_locks_lower_in(6,20) <= s_locks_lower_out(7,20);

		normal_cell_6_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,21),
			fetch              => s_fetch(6,21),
			data_in            => s_data_in(6,21),
			data_out           => s_data_out(6,21),
			out1               => s_out1(6,21),
			out2               => s_out2(6,21),
			lock_lower_row_out => s_locks_lower_out(6,21),
			lock_lower_row_in  => s_locks_lower_in(6,21),
			in1                => s_in1(6,21),
			in2                => s_in2(6,21),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(21)
		);
	s_in1(6,21)            <= s_out1(7,21);
	s_in2(6,21)            <= s_out2(7,22);
	s_locks_lower_in(6,21) <= s_locks_lower_out(7,21);

		normal_cell_6_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,22),
			fetch              => s_fetch(6,22),
			data_in            => s_data_in(6,22),
			data_out           => s_data_out(6,22),
			out1               => s_out1(6,22),
			out2               => s_out2(6,22),
			lock_lower_row_out => s_locks_lower_out(6,22),
			lock_lower_row_in  => s_locks_lower_in(6,22),
			in1                => s_in1(6,22),
			in2                => s_in2(6,22),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(22)
		);
	s_in1(6,22)            <= s_out1(7,22);
	s_in2(6,22)            <= s_out2(7,23);
	s_locks_lower_in(6,22) <= s_locks_lower_out(7,22);

		normal_cell_6_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,23),
			fetch              => s_fetch(6,23),
			data_in            => s_data_in(6,23),
			data_out           => s_data_out(6,23),
			out1               => s_out1(6,23),
			out2               => s_out2(6,23),
			lock_lower_row_out => s_locks_lower_out(6,23),
			lock_lower_row_in  => s_locks_lower_in(6,23),
			in1                => s_in1(6,23),
			in2                => s_in2(6,23),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(23)
		);
	s_in1(6,23)            <= s_out1(7,23);
	s_in2(6,23)            <= s_out2(7,24);
	s_locks_lower_in(6,23) <= s_locks_lower_out(7,23);

		normal_cell_6_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,24),
			fetch              => s_fetch(6,24),
			data_in            => s_data_in(6,24),
			data_out           => s_data_out(6,24),
			out1               => s_out1(6,24),
			out2               => s_out2(6,24),
			lock_lower_row_out => s_locks_lower_out(6,24),
			lock_lower_row_in  => s_locks_lower_in(6,24),
			in1                => s_in1(6,24),
			in2                => s_in2(6,24),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(24)
		);
	s_in1(6,24)            <= s_out1(7,24);
	s_in2(6,24)            <= s_out2(7,25);
	s_locks_lower_in(6,24) <= s_locks_lower_out(7,24);

		normal_cell_6_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,25),
			fetch              => s_fetch(6,25),
			data_in            => s_data_in(6,25),
			data_out           => s_data_out(6,25),
			out1               => s_out1(6,25),
			out2               => s_out2(6,25),
			lock_lower_row_out => s_locks_lower_out(6,25),
			lock_lower_row_in  => s_locks_lower_in(6,25),
			in1                => s_in1(6,25),
			in2                => s_in2(6,25),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(25)
		);
	s_in1(6,25)            <= s_out1(7,25);
	s_in2(6,25)            <= s_out2(7,26);
	s_locks_lower_in(6,25) <= s_locks_lower_out(7,25);

		normal_cell_6_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,26),
			fetch              => s_fetch(6,26),
			data_in            => s_data_in(6,26),
			data_out           => s_data_out(6,26),
			out1               => s_out1(6,26),
			out2               => s_out2(6,26),
			lock_lower_row_out => s_locks_lower_out(6,26),
			lock_lower_row_in  => s_locks_lower_in(6,26),
			in1                => s_in1(6,26),
			in2                => s_in2(6,26),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(26)
		);
	s_in1(6,26)            <= s_out1(7,26);
	s_in2(6,26)            <= s_out2(7,27);
	s_locks_lower_in(6,26) <= s_locks_lower_out(7,26);

		normal_cell_6_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,27),
			fetch              => s_fetch(6,27),
			data_in            => s_data_in(6,27),
			data_out           => s_data_out(6,27),
			out1               => s_out1(6,27),
			out2               => s_out2(6,27),
			lock_lower_row_out => s_locks_lower_out(6,27),
			lock_lower_row_in  => s_locks_lower_in(6,27),
			in1                => s_in1(6,27),
			in2                => s_in2(6,27),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(27)
		);
	s_in1(6,27)            <= s_out1(7,27);
	s_in2(6,27)            <= s_out2(7,28);
	s_locks_lower_in(6,27) <= s_locks_lower_out(7,27);

		normal_cell_6_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,28),
			fetch              => s_fetch(6,28),
			data_in            => s_data_in(6,28),
			data_out           => s_data_out(6,28),
			out1               => s_out1(6,28),
			out2               => s_out2(6,28),
			lock_lower_row_out => s_locks_lower_out(6,28),
			lock_lower_row_in  => s_locks_lower_in(6,28),
			in1                => s_in1(6,28),
			in2                => s_in2(6,28),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(28)
		);
	s_in1(6,28)            <= s_out1(7,28);
	s_in2(6,28)            <= s_out2(7,29);
	s_locks_lower_in(6,28) <= s_locks_lower_out(7,28);

		normal_cell_6_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,29),
			fetch              => s_fetch(6,29),
			data_in            => s_data_in(6,29),
			data_out           => s_data_out(6,29),
			out1               => s_out1(6,29),
			out2               => s_out2(6,29),
			lock_lower_row_out => s_locks_lower_out(6,29),
			lock_lower_row_in  => s_locks_lower_in(6,29),
			in1                => s_in1(6,29),
			in2                => s_in2(6,29),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(29)
		);
	s_in1(6,29)            <= s_out1(7,29);
	s_in2(6,29)            <= s_out2(7,30);
	s_locks_lower_in(6,29) <= s_locks_lower_out(7,29);

		normal_cell_6_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,30),
			fetch              => s_fetch(6,30),
			data_in            => s_data_in(6,30),
			data_out           => s_data_out(6,30),
			out1               => s_out1(6,30),
			out2               => s_out2(6,30),
			lock_lower_row_out => s_locks_lower_out(6,30),
			lock_lower_row_in  => s_locks_lower_in(6,30),
			in1                => s_in1(6,30),
			in2                => s_in2(6,30),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(30)
		);
	s_in1(6,30)            <= s_out1(7,30);
	s_in2(6,30)            <= s_out2(7,31);
	s_locks_lower_in(6,30) <= s_locks_lower_out(7,30);

		normal_cell_6_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,31),
			fetch              => s_fetch(6,31),
			data_in            => s_data_in(6,31),
			data_out           => s_data_out(6,31),
			out1               => s_out1(6,31),
			out2               => s_out2(6,31),
			lock_lower_row_out => s_locks_lower_out(6,31),
			lock_lower_row_in  => s_locks_lower_in(6,31),
			in1                => s_in1(6,31),
			in2                => s_in2(6,31),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(31)
		);
	s_in1(6,31)            <= s_out1(7,31);
	s_in2(6,31)            <= s_out2(7,32);
	s_locks_lower_in(6,31) <= s_locks_lower_out(7,31);

		normal_cell_6_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,32),
			fetch              => s_fetch(6,32),
			data_in            => s_data_in(6,32),
			data_out           => s_data_out(6,32),
			out1               => s_out1(6,32),
			out2               => s_out2(6,32),
			lock_lower_row_out => s_locks_lower_out(6,32),
			lock_lower_row_in  => s_locks_lower_in(6,32),
			in1                => s_in1(6,32),
			in2                => s_in2(6,32),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(32)
		);
	s_in1(6,32)            <= s_out1(7,32);
	s_in2(6,32)            <= s_out2(7,33);
	s_locks_lower_in(6,32) <= s_locks_lower_out(7,32);

		normal_cell_6_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,33),
			fetch              => s_fetch(6,33),
			data_in            => s_data_in(6,33),
			data_out           => s_data_out(6,33),
			out1               => s_out1(6,33),
			out2               => s_out2(6,33),
			lock_lower_row_out => s_locks_lower_out(6,33),
			lock_lower_row_in  => s_locks_lower_in(6,33),
			in1                => s_in1(6,33),
			in2                => s_in2(6,33),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(33)
		);
	s_in1(6,33)            <= s_out1(7,33);
	s_in2(6,33)            <= s_out2(7,34);
	s_locks_lower_in(6,33) <= s_locks_lower_out(7,33);

		normal_cell_6_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,34),
			fetch              => s_fetch(6,34),
			data_in            => s_data_in(6,34),
			data_out           => s_data_out(6,34),
			out1               => s_out1(6,34),
			out2               => s_out2(6,34),
			lock_lower_row_out => s_locks_lower_out(6,34),
			lock_lower_row_in  => s_locks_lower_in(6,34),
			in1                => s_in1(6,34),
			in2                => s_in2(6,34),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(34)
		);
	s_in1(6,34)            <= s_out1(7,34);
	s_in2(6,34)            <= s_out2(7,35);
	s_locks_lower_in(6,34) <= s_locks_lower_out(7,34);

		normal_cell_6_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,35),
			fetch              => s_fetch(6,35),
			data_in            => s_data_in(6,35),
			data_out           => s_data_out(6,35),
			out1               => s_out1(6,35),
			out2               => s_out2(6,35),
			lock_lower_row_out => s_locks_lower_out(6,35),
			lock_lower_row_in  => s_locks_lower_in(6,35),
			in1                => s_in1(6,35),
			in2                => s_in2(6,35),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(35)
		);
	s_in1(6,35)            <= s_out1(7,35);
	s_in2(6,35)            <= s_out2(7,36);
	s_locks_lower_in(6,35) <= s_locks_lower_out(7,35);

		normal_cell_6_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,36),
			fetch              => s_fetch(6,36),
			data_in            => s_data_in(6,36),
			data_out           => s_data_out(6,36),
			out1               => s_out1(6,36),
			out2               => s_out2(6,36),
			lock_lower_row_out => s_locks_lower_out(6,36),
			lock_lower_row_in  => s_locks_lower_in(6,36),
			in1                => s_in1(6,36),
			in2                => s_in2(6,36),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(36)
		);
	s_in1(6,36)            <= s_out1(7,36);
	s_in2(6,36)            <= s_out2(7,37);
	s_locks_lower_in(6,36) <= s_locks_lower_out(7,36);

		normal_cell_6_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,37),
			fetch              => s_fetch(6,37),
			data_in            => s_data_in(6,37),
			data_out           => s_data_out(6,37),
			out1               => s_out1(6,37),
			out2               => s_out2(6,37),
			lock_lower_row_out => s_locks_lower_out(6,37),
			lock_lower_row_in  => s_locks_lower_in(6,37),
			in1                => s_in1(6,37),
			in2                => s_in2(6,37),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(37)
		);
	s_in1(6,37)            <= s_out1(7,37);
	s_in2(6,37)            <= s_out2(7,38);
	s_locks_lower_in(6,37) <= s_locks_lower_out(7,37);

		normal_cell_6_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,38),
			fetch              => s_fetch(6,38),
			data_in            => s_data_in(6,38),
			data_out           => s_data_out(6,38),
			out1               => s_out1(6,38),
			out2               => s_out2(6,38),
			lock_lower_row_out => s_locks_lower_out(6,38),
			lock_lower_row_in  => s_locks_lower_in(6,38),
			in1                => s_in1(6,38),
			in2                => s_in2(6,38),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(38)
		);
	s_in1(6,38)            <= s_out1(7,38);
	s_in2(6,38)            <= s_out2(7,39);
	s_locks_lower_in(6,38) <= s_locks_lower_out(7,38);

		normal_cell_6_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,39),
			fetch              => s_fetch(6,39),
			data_in            => s_data_in(6,39),
			data_out           => s_data_out(6,39),
			out1               => s_out1(6,39),
			out2               => s_out2(6,39),
			lock_lower_row_out => s_locks_lower_out(6,39),
			lock_lower_row_in  => s_locks_lower_in(6,39),
			in1                => s_in1(6,39),
			in2                => s_in2(6,39),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(39)
		);
	s_in1(6,39)            <= s_out1(7,39);
	s_in2(6,39)            <= s_out2(7,40);
	s_locks_lower_in(6,39) <= s_locks_lower_out(7,39);

		normal_cell_6_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,40),
			fetch              => s_fetch(6,40),
			data_in            => s_data_in(6,40),
			data_out           => s_data_out(6,40),
			out1               => s_out1(6,40),
			out2               => s_out2(6,40),
			lock_lower_row_out => s_locks_lower_out(6,40),
			lock_lower_row_in  => s_locks_lower_in(6,40),
			in1                => s_in1(6,40),
			in2                => s_in2(6,40),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(40)
		);
	s_in1(6,40)            <= s_out1(7,40);
	s_in2(6,40)            <= s_out2(7,41);
	s_locks_lower_in(6,40) <= s_locks_lower_out(7,40);

		normal_cell_6_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,41),
			fetch              => s_fetch(6,41),
			data_in            => s_data_in(6,41),
			data_out           => s_data_out(6,41),
			out1               => s_out1(6,41),
			out2               => s_out2(6,41),
			lock_lower_row_out => s_locks_lower_out(6,41),
			lock_lower_row_in  => s_locks_lower_in(6,41),
			in1                => s_in1(6,41),
			in2                => s_in2(6,41),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(41)
		);
	s_in1(6,41)            <= s_out1(7,41);
	s_in2(6,41)            <= s_out2(7,42);
	s_locks_lower_in(6,41) <= s_locks_lower_out(7,41);

		normal_cell_6_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,42),
			fetch              => s_fetch(6,42),
			data_in            => s_data_in(6,42),
			data_out           => s_data_out(6,42),
			out1               => s_out1(6,42),
			out2               => s_out2(6,42),
			lock_lower_row_out => s_locks_lower_out(6,42),
			lock_lower_row_in  => s_locks_lower_in(6,42),
			in1                => s_in1(6,42),
			in2                => s_in2(6,42),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(42)
		);
	s_in1(6,42)            <= s_out1(7,42);
	s_in2(6,42)            <= s_out2(7,43);
	s_locks_lower_in(6,42) <= s_locks_lower_out(7,42);

		normal_cell_6_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,43),
			fetch              => s_fetch(6,43),
			data_in            => s_data_in(6,43),
			data_out           => s_data_out(6,43),
			out1               => s_out1(6,43),
			out2               => s_out2(6,43),
			lock_lower_row_out => s_locks_lower_out(6,43),
			lock_lower_row_in  => s_locks_lower_in(6,43),
			in1                => s_in1(6,43),
			in2                => s_in2(6,43),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(43)
		);
	s_in1(6,43)            <= s_out1(7,43);
	s_in2(6,43)            <= s_out2(7,44);
	s_locks_lower_in(6,43) <= s_locks_lower_out(7,43);

		normal_cell_6_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,44),
			fetch              => s_fetch(6,44),
			data_in            => s_data_in(6,44),
			data_out           => s_data_out(6,44),
			out1               => s_out1(6,44),
			out2               => s_out2(6,44),
			lock_lower_row_out => s_locks_lower_out(6,44),
			lock_lower_row_in  => s_locks_lower_in(6,44),
			in1                => s_in1(6,44),
			in2                => s_in2(6,44),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(44)
		);
	s_in1(6,44)            <= s_out1(7,44);
	s_in2(6,44)            <= s_out2(7,45);
	s_locks_lower_in(6,44) <= s_locks_lower_out(7,44);

		normal_cell_6_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,45),
			fetch              => s_fetch(6,45),
			data_in            => s_data_in(6,45),
			data_out           => s_data_out(6,45),
			out1               => s_out1(6,45),
			out2               => s_out2(6,45),
			lock_lower_row_out => s_locks_lower_out(6,45),
			lock_lower_row_in  => s_locks_lower_in(6,45),
			in1                => s_in1(6,45),
			in2                => s_in2(6,45),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(45)
		);
	s_in1(6,45)            <= s_out1(7,45);
	s_in2(6,45)            <= s_out2(7,46);
	s_locks_lower_in(6,45) <= s_locks_lower_out(7,45);

		normal_cell_6_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,46),
			fetch              => s_fetch(6,46),
			data_in            => s_data_in(6,46),
			data_out           => s_data_out(6,46),
			out1               => s_out1(6,46),
			out2               => s_out2(6,46),
			lock_lower_row_out => s_locks_lower_out(6,46),
			lock_lower_row_in  => s_locks_lower_in(6,46),
			in1                => s_in1(6,46),
			in2                => s_in2(6,46),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(46)
		);
	s_in1(6,46)            <= s_out1(7,46);
	s_in2(6,46)            <= s_out2(7,47);
	s_locks_lower_in(6,46) <= s_locks_lower_out(7,46);

		normal_cell_6_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,47),
			fetch              => s_fetch(6,47),
			data_in            => s_data_in(6,47),
			data_out           => s_data_out(6,47),
			out1               => s_out1(6,47),
			out2               => s_out2(6,47),
			lock_lower_row_out => s_locks_lower_out(6,47),
			lock_lower_row_in  => s_locks_lower_in(6,47),
			in1                => s_in1(6,47),
			in2                => s_in2(6,47),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(47)
		);
	s_in1(6,47)            <= s_out1(7,47);
	s_in2(6,47)            <= s_out2(7,48);
	s_locks_lower_in(6,47) <= s_locks_lower_out(7,47);

		normal_cell_6_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,48),
			fetch              => s_fetch(6,48),
			data_in            => s_data_in(6,48),
			data_out           => s_data_out(6,48),
			out1               => s_out1(6,48),
			out2               => s_out2(6,48),
			lock_lower_row_out => s_locks_lower_out(6,48),
			lock_lower_row_in  => s_locks_lower_in(6,48),
			in1                => s_in1(6,48),
			in2                => s_in2(6,48),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(48)
		);
	s_in1(6,48)            <= s_out1(7,48);
	s_in2(6,48)            <= s_out2(7,49);
	s_locks_lower_in(6,48) <= s_locks_lower_out(7,48);

		normal_cell_6_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,49),
			fetch              => s_fetch(6,49),
			data_in            => s_data_in(6,49),
			data_out           => s_data_out(6,49),
			out1               => s_out1(6,49),
			out2               => s_out2(6,49),
			lock_lower_row_out => s_locks_lower_out(6,49),
			lock_lower_row_in  => s_locks_lower_in(6,49),
			in1                => s_in1(6,49),
			in2                => s_in2(6,49),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(49)
		);
	s_in1(6,49)            <= s_out1(7,49);
	s_in2(6,49)            <= s_out2(7,50);
	s_locks_lower_in(6,49) <= s_locks_lower_out(7,49);

		normal_cell_6_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,50),
			fetch              => s_fetch(6,50),
			data_in            => s_data_in(6,50),
			data_out           => s_data_out(6,50),
			out1               => s_out1(6,50),
			out2               => s_out2(6,50),
			lock_lower_row_out => s_locks_lower_out(6,50),
			lock_lower_row_in  => s_locks_lower_in(6,50),
			in1                => s_in1(6,50),
			in2                => s_in2(6,50),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(50)
		);
	s_in1(6,50)            <= s_out1(7,50);
	s_in2(6,50)            <= s_out2(7,51);
	s_locks_lower_in(6,50) <= s_locks_lower_out(7,50);

		normal_cell_6_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,51),
			fetch              => s_fetch(6,51),
			data_in            => s_data_in(6,51),
			data_out           => s_data_out(6,51),
			out1               => s_out1(6,51),
			out2               => s_out2(6,51),
			lock_lower_row_out => s_locks_lower_out(6,51),
			lock_lower_row_in  => s_locks_lower_in(6,51),
			in1                => s_in1(6,51),
			in2                => s_in2(6,51),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(51)
		);
	s_in1(6,51)            <= s_out1(7,51);
	s_in2(6,51)            <= s_out2(7,52);
	s_locks_lower_in(6,51) <= s_locks_lower_out(7,51);

		normal_cell_6_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,52),
			fetch              => s_fetch(6,52),
			data_in            => s_data_in(6,52),
			data_out           => s_data_out(6,52),
			out1               => s_out1(6,52),
			out2               => s_out2(6,52),
			lock_lower_row_out => s_locks_lower_out(6,52),
			lock_lower_row_in  => s_locks_lower_in(6,52),
			in1                => s_in1(6,52),
			in2                => s_in2(6,52),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(52)
		);
	s_in1(6,52)            <= s_out1(7,52);
	s_in2(6,52)            <= s_out2(7,53);
	s_locks_lower_in(6,52) <= s_locks_lower_out(7,52);

		normal_cell_6_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,53),
			fetch              => s_fetch(6,53),
			data_in            => s_data_in(6,53),
			data_out           => s_data_out(6,53),
			out1               => s_out1(6,53),
			out2               => s_out2(6,53),
			lock_lower_row_out => s_locks_lower_out(6,53),
			lock_lower_row_in  => s_locks_lower_in(6,53),
			in1                => s_in1(6,53),
			in2                => s_in2(6,53),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(53)
		);
	s_in1(6,53)            <= s_out1(7,53);
	s_in2(6,53)            <= s_out2(7,54);
	s_locks_lower_in(6,53) <= s_locks_lower_out(7,53);

		normal_cell_6_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,54),
			fetch              => s_fetch(6,54),
			data_in            => s_data_in(6,54),
			data_out           => s_data_out(6,54),
			out1               => s_out1(6,54),
			out2               => s_out2(6,54),
			lock_lower_row_out => s_locks_lower_out(6,54),
			lock_lower_row_in  => s_locks_lower_in(6,54),
			in1                => s_in1(6,54),
			in2                => s_in2(6,54),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(54)
		);
	s_in1(6,54)            <= s_out1(7,54);
	s_in2(6,54)            <= s_out2(7,55);
	s_locks_lower_in(6,54) <= s_locks_lower_out(7,54);

		normal_cell_6_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,55),
			fetch              => s_fetch(6,55),
			data_in            => s_data_in(6,55),
			data_out           => s_data_out(6,55),
			out1               => s_out1(6,55),
			out2               => s_out2(6,55),
			lock_lower_row_out => s_locks_lower_out(6,55),
			lock_lower_row_in  => s_locks_lower_in(6,55),
			in1                => s_in1(6,55),
			in2                => s_in2(6,55),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(55)
		);
	s_in1(6,55)            <= s_out1(7,55);
	s_in2(6,55)            <= s_out2(7,56);
	s_locks_lower_in(6,55) <= s_locks_lower_out(7,55);

		normal_cell_6_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,56),
			fetch              => s_fetch(6,56),
			data_in            => s_data_in(6,56),
			data_out           => s_data_out(6,56),
			out1               => s_out1(6,56),
			out2               => s_out2(6,56),
			lock_lower_row_out => s_locks_lower_out(6,56),
			lock_lower_row_in  => s_locks_lower_in(6,56),
			in1                => s_in1(6,56),
			in2                => s_in2(6,56),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(56)
		);
	s_in1(6,56)            <= s_out1(7,56);
	s_in2(6,56)            <= s_out2(7,57);
	s_locks_lower_in(6,56) <= s_locks_lower_out(7,56);

		normal_cell_6_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,57),
			fetch              => s_fetch(6,57),
			data_in            => s_data_in(6,57),
			data_out           => s_data_out(6,57),
			out1               => s_out1(6,57),
			out2               => s_out2(6,57),
			lock_lower_row_out => s_locks_lower_out(6,57),
			lock_lower_row_in  => s_locks_lower_in(6,57),
			in1                => s_in1(6,57),
			in2                => s_in2(6,57),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(57)
		);
	s_in1(6,57)            <= s_out1(7,57);
	s_in2(6,57)            <= s_out2(7,58);
	s_locks_lower_in(6,57) <= s_locks_lower_out(7,57);

		normal_cell_6_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,58),
			fetch              => s_fetch(6,58),
			data_in            => s_data_in(6,58),
			data_out           => s_data_out(6,58),
			out1               => s_out1(6,58),
			out2               => s_out2(6,58),
			lock_lower_row_out => s_locks_lower_out(6,58),
			lock_lower_row_in  => s_locks_lower_in(6,58),
			in1                => s_in1(6,58),
			in2                => s_in2(6,58),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(58)
		);
	s_in1(6,58)            <= s_out1(7,58);
	s_in2(6,58)            <= s_out2(7,59);
	s_locks_lower_in(6,58) <= s_locks_lower_out(7,58);

		normal_cell_6_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,59),
			fetch              => s_fetch(6,59),
			data_in            => s_data_in(6,59),
			data_out           => s_data_out(6,59),
			out1               => s_out1(6,59),
			out2               => s_out2(6,59),
			lock_lower_row_out => s_locks_lower_out(6,59),
			lock_lower_row_in  => s_locks_lower_in(6,59),
			in1                => s_in1(6,59),
			in2                => s_in2(6,59),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(59)
		);
	s_in1(6,59)            <= s_out1(7,59);
	s_in2(6,59)            <= s_out2(7,60);
	s_locks_lower_in(6,59) <= s_locks_lower_out(7,59);

		last_col_cell_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(6,60),
			fetch              => s_fetch(6,60),
			data_in            => s_data_in(6,60),
			data_out           => s_data_out(6,60),
			out1               => s_out1(6,60),
			out2               => s_out2(6,60),
			lock_lower_row_out => s_locks_lower_out(6,60),
			lock_lower_row_in  => s_locks_lower_in(6,60),
			in1                => s_in1(6,60),
			in2                => (others => '0'),
			lock_row           => s_locks(6),
			piv_found          => s_piv_found,
			row_data           => s_row_data(6),
			col_data           => s_col_data(60)
		);
	s_in1(6,60)            <= s_out1(7,60);
	s_locks_lower_in(6,60) <= s_locks_lower_out(7,60);

		normal_cell_7_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,1),
			fetch              => s_fetch(7,1),
			data_in            => s_data_in(7,1),
			data_out           => s_data_out(7,1),
			out1               => s_out1(7,1),
			out2               => s_out2(7,1),
			lock_lower_row_out => s_locks_lower_out(7,1),
			lock_lower_row_in  => s_locks_lower_in(7,1),
			in1                => s_in1(7,1),
			in2                => s_in2(7,1),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(1)
		);
	s_in1(7,1)            <= s_out1(8,1);
	s_in2(7,1)            <= s_out2(8,2);
	s_locks_lower_in(7,1) <= s_locks_lower_out(8,1);

		normal_cell_7_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,2),
			fetch              => s_fetch(7,2),
			data_in            => s_data_in(7,2),
			data_out           => s_data_out(7,2),
			out1               => s_out1(7,2),
			out2               => s_out2(7,2),
			lock_lower_row_out => s_locks_lower_out(7,2),
			lock_lower_row_in  => s_locks_lower_in(7,2),
			in1                => s_in1(7,2),
			in2                => s_in2(7,2),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(2)
		);
	s_in1(7,2)            <= s_out1(8,2);
	s_in2(7,2)            <= s_out2(8,3);
	s_locks_lower_in(7,2) <= s_locks_lower_out(8,2);

		normal_cell_7_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,3),
			fetch              => s_fetch(7,3),
			data_in            => s_data_in(7,3),
			data_out           => s_data_out(7,3),
			out1               => s_out1(7,3),
			out2               => s_out2(7,3),
			lock_lower_row_out => s_locks_lower_out(7,3),
			lock_lower_row_in  => s_locks_lower_in(7,3),
			in1                => s_in1(7,3),
			in2                => s_in2(7,3),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(3)
		);
	s_in1(7,3)            <= s_out1(8,3);
	s_in2(7,3)            <= s_out2(8,4);
	s_locks_lower_in(7,3) <= s_locks_lower_out(8,3);

		normal_cell_7_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,4),
			fetch              => s_fetch(7,4),
			data_in            => s_data_in(7,4),
			data_out           => s_data_out(7,4),
			out1               => s_out1(7,4),
			out2               => s_out2(7,4),
			lock_lower_row_out => s_locks_lower_out(7,4),
			lock_lower_row_in  => s_locks_lower_in(7,4),
			in1                => s_in1(7,4),
			in2                => s_in2(7,4),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(4)
		);
	s_in1(7,4)            <= s_out1(8,4);
	s_in2(7,4)            <= s_out2(8,5);
	s_locks_lower_in(7,4) <= s_locks_lower_out(8,4);

		normal_cell_7_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,5),
			fetch              => s_fetch(7,5),
			data_in            => s_data_in(7,5),
			data_out           => s_data_out(7,5),
			out1               => s_out1(7,5),
			out2               => s_out2(7,5),
			lock_lower_row_out => s_locks_lower_out(7,5),
			lock_lower_row_in  => s_locks_lower_in(7,5),
			in1                => s_in1(7,5),
			in2                => s_in2(7,5),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(5)
		);
	s_in1(7,5)            <= s_out1(8,5);
	s_in2(7,5)            <= s_out2(8,6);
	s_locks_lower_in(7,5) <= s_locks_lower_out(8,5);

		normal_cell_7_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,6),
			fetch              => s_fetch(7,6),
			data_in            => s_data_in(7,6),
			data_out           => s_data_out(7,6),
			out1               => s_out1(7,6),
			out2               => s_out2(7,6),
			lock_lower_row_out => s_locks_lower_out(7,6),
			lock_lower_row_in  => s_locks_lower_in(7,6),
			in1                => s_in1(7,6),
			in2                => s_in2(7,6),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(6)
		);
	s_in1(7,6)            <= s_out1(8,6);
	s_in2(7,6)            <= s_out2(8,7);
	s_locks_lower_in(7,6) <= s_locks_lower_out(8,6);

		normal_cell_7_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,7),
			fetch              => s_fetch(7,7),
			data_in            => s_data_in(7,7),
			data_out           => s_data_out(7,7),
			out1               => s_out1(7,7),
			out2               => s_out2(7,7),
			lock_lower_row_out => s_locks_lower_out(7,7),
			lock_lower_row_in  => s_locks_lower_in(7,7),
			in1                => s_in1(7,7),
			in2                => s_in2(7,7),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(7)
		);
	s_in1(7,7)            <= s_out1(8,7);
	s_in2(7,7)            <= s_out2(8,8);
	s_locks_lower_in(7,7) <= s_locks_lower_out(8,7);

		normal_cell_7_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,8),
			fetch              => s_fetch(7,8),
			data_in            => s_data_in(7,8),
			data_out           => s_data_out(7,8),
			out1               => s_out1(7,8),
			out2               => s_out2(7,8),
			lock_lower_row_out => s_locks_lower_out(7,8),
			lock_lower_row_in  => s_locks_lower_in(7,8),
			in1                => s_in1(7,8),
			in2                => s_in2(7,8),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(8)
		);
	s_in1(7,8)            <= s_out1(8,8);
	s_in2(7,8)            <= s_out2(8,9);
	s_locks_lower_in(7,8) <= s_locks_lower_out(8,8);

		normal_cell_7_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,9),
			fetch              => s_fetch(7,9),
			data_in            => s_data_in(7,9),
			data_out           => s_data_out(7,9),
			out1               => s_out1(7,9),
			out2               => s_out2(7,9),
			lock_lower_row_out => s_locks_lower_out(7,9),
			lock_lower_row_in  => s_locks_lower_in(7,9),
			in1                => s_in1(7,9),
			in2                => s_in2(7,9),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(9)
		);
	s_in1(7,9)            <= s_out1(8,9);
	s_in2(7,9)            <= s_out2(8,10);
	s_locks_lower_in(7,9) <= s_locks_lower_out(8,9);

		normal_cell_7_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,10),
			fetch              => s_fetch(7,10),
			data_in            => s_data_in(7,10),
			data_out           => s_data_out(7,10),
			out1               => s_out1(7,10),
			out2               => s_out2(7,10),
			lock_lower_row_out => s_locks_lower_out(7,10),
			lock_lower_row_in  => s_locks_lower_in(7,10),
			in1                => s_in1(7,10),
			in2                => s_in2(7,10),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(10)
		);
	s_in1(7,10)            <= s_out1(8,10);
	s_in2(7,10)            <= s_out2(8,11);
	s_locks_lower_in(7,10) <= s_locks_lower_out(8,10);

		normal_cell_7_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,11),
			fetch              => s_fetch(7,11),
			data_in            => s_data_in(7,11),
			data_out           => s_data_out(7,11),
			out1               => s_out1(7,11),
			out2               => s_out2(7,11),
			lock_lower_row_out => s_locks_lower_out(7,11),
			lock_lower_row_in  => s_locks_lower_in(7,11),
			in1                => s_in1(7,11),
			in2                => s_in2(7,11),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(11)
		);
	s_in1(7,11)            <= s_out1(8,11);
	s_in2(7,11)            <= s_out2(8,12);
	s_locks_lower_in(7,11) <= s_locks_lower_out(8,11);

		normal_cell_7_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,12),
			fetch              => s_fetch(7,12),
			data_in            => s_data_in(7,12),
			data_out           => s_data_out(7,12),
			out1               => s_out1(7,12),
			out2               => s_out2(7,12),
			lock_lower_row_out => s_locks_lower_out(7,12),
			lock_lower_row_in  => s_locks_lower_in(7,12),
			in1                => s_in1(7,12),
			in2                => s_in2(7,12),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(12)
		);
	s_in1(7,12)            <= s_out1(8,12);
	s_in2(7,12)            <= s_out2(8,13);
	s_locks_lower_in(7,12) <= s_locks_lower_out(8,12);

		normal_cell_7_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,13),
			fetch              => s_fetch(7,13),
			data_in            => s_data_in(7,13),
			data_out           => s_data_out(7,13),
			out1               => s_out1(7,13),
			out2               => s_out2(7,13),
			lock_lower_row_out => s_locks_lower_out(7,13),
			lock_lower_row_in  => s_locks_lower_in(7,13),
			in1                => s_in1(7,13),
			in2                => s_in2(7,13),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(13)
		);
	s_in1(7,13)            <= s_out1(8,13);
	s_in2(7,13)            <= s_out2(8,14);
	s_locks_lower_in(7,13) <= s_locks_lower_out(8,13);

		normal_cell_7_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,14),
			fetch              => s_fetch(7,14),
			data_in            => s_data_in(7,14),
			data_out           => s_data_out(7,14),
			out1               => s_out1(7,14),
			out2               => s_out2(7,14),
			lock_lower_row_out => s_locks_lower_out(7,14),
			lock_lower_row_in  => s_locks_lower_in(7,14),
			in1                => s_in1(7,14),
			in2                => s_in2(7,14),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(14)
		);
	s_in1(7,14)            <= s_out1(8,14);
	s_in2(7,14)            <= s_out2(8,15);
	s_locks_lower_in(7,14) <= s_locks_lower_out(8,14);

		normal_cell_7_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,15),
			fetch              => s_fetch(7,15),
			data_in            => s_data_in(7,15),
			data_out           => s_data_out(7,15),
			out1               => s_out1(7,15),
			out2               => s_out2(7,15),
			lock_lower_row_out => s_locks_lower_out(7,15),
			lock_lower_row_in  => s_locks_lower_in(7,15),
			in1                => s_in1(7,15),
			in2                => s_in2(7,15),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(15)
		);
	s_in1(7,15)            <= s_out1(8,15);
	s_in2(7,15)            <= s_out2(8,16);
	s_locks_lower_in(7,15) <= s_locks_lower_out(8,15);

		normal_cell_7_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,16),
			fetch              => s_fetch(7,16),
			data_in            => s_data_in(7,16),
			data_out           => s_data_out(7,16),
			out1               => s_out1(7,16),
			out2               => s_out2(7,16),
			lock_lower_row_out => s_locks_lower_out(7,16),
			lock_lower_row_in  => s_locks_lower_in(7,16),
			in1                => s_in1(7,16),
			in2                => s_in2(7,16),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(16)
		);
	s_in1(7,16)            <= s_out1(8,16);
	s_in2(7,16)            <= s_out2(8,17);
	s_locks_lower_in(7,16) <= s_locks_lower_out(8,16);

		normal_cell_7_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,17),
			fetch              => s_fetch(7,17),
			data_in            => s_data_in(7,17),
			data_out           => s_data_out(7,17),
			out1               => s_out1(7,17),
			out2               => s_out2(7,17),
			lock_lower_row_out => s_locks_lower_out(7,17),
			lock_lower_row_in  => s_locks_lower_in(7,17),
			in1                => s_in1(7,17),
			in2                => s_in2(7,17),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(17)
		);
	s_in1(7,17)            <= s_out1(8,17);
	s_in2(7,17)            <= s_out2(8,18);
	s_locks_lower_in(7,17) <= s_locks_lower_out(8,17);

		normal_cell_7_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,18),
			fetch              => s_fetch(7,18),
			data_in            => s_data_in(7,18),
			data_out           => s_data_out(7,18),
			out1               => s_out1(7,18),
			out2               => s_out2(7,18),
			lock_lower_row_out => s_locks_lower_out(7,18),
			lock_lower_row_in  => s_locks_lower_in(7,18),
			in1                => s_in1(7,18),
			in2                => s_in2(7,18),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(18)
		);
	s_in1(7,18)            <= s_out1(8,18);
	s_in2(7,18)            <= s_out2(8,19);
	s_locks_lower_in(7,18) <= s_locks_lower_out(8,18);

		normal_cell_7_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,19),
			fetch              => s_fetch(7,19),
			data_in            => s_data_in(7,19),
			data_out           => s_data_out(7,19),
			out1               => s_out1(7,19),
			out2               => s_out2(7,19),
			lock_lower_row_out => s_locks_lower_out(7,19),
			lock_lower_row_in  => s_locks_lower_in(7,19),
			in1                => s_in1(7,19),
			in2                => s_in2(7,19),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(19)
		);
	s_in1(7,19)            <= s_out1(8,19);
	s_in2(7,19)            <= s_out2(8,20);
	s_locks_lower_in(7,19) <= s_locks_lower_out(8,19);

		normal_cell_7_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,20),
			fetch              => s_fetch(7,20),
			data_in            => s_data_in(7,20),
			data_out           => s_data_out(7,20),
			out1               => s_out1(7,20),
			out2               => s_out2(7,20),
			lock_lower_row_out => s_locks_lower_out(7,20),
			lock_lower_row_in  => s_locks_lower_in(7,20),
			in1                => s_in1(7,20),
			in2                => s_in2(7,20),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(20)
		);
	s_in1(7,20)            <= s_out1(8,20);
	s_in2(7,20)            <= s_out2(8,21);
	s_locks_lower_in(7,20) <= s_locks_lower_out(8,20);

		normal_cell_7_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,21),
			fetch              => s_fetch(7,21),
			data_in            => s_data_in(7,21),
			data_out           => s_data_out(7,21),
			out1               => s_out1(7,21),
			out2               => s_out2(7,21),
			lock_lower_row_out => s_locks_lower_out(7,21),
			lock_lower_row_in  => s_locks_lower_in(7,21),
			in1                => s_in1(7,21),
			in2                => s_in2(7,21),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(21)
		);
	s_in1(7,21)            <= s_out1(8,21);
	s_in2(7,21)            <= s_out2(8,22);
	s_locks_lower_in(7,21) <= s_locks_lower_out(8,21);

		normal_cell_7_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,22),
			fetch              => s_fetch(7,22),
			data_in            => s_data_in(7,22),
			data_out           => s_data_out(7,22),
			out1               => s_out1(7,22),
			out2               => s_out2(7,22),
			lock_lower_row_out => s_locks_lower_out(7,22),
			lock_lower_row_in  => s_locks_lower_in(7,22),
			in1                => s_in1(7,22),
			in2                => s_in2(7,22),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(22)
		);
	s_in1(7,22)            <= s_out1(8,22);
	s_in2(7,22)            <= s_out2(8,23);
	s_locks_lower_in(7,22) <= s_locks_lower_out(8,22);

		normal_cell_7_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,23),
			fetch              => s_fetch(7,23),
			data_in            => s_data_in(7,23),
			data_out           => s_data_out(7,23),
			out1               => s_out1(7,23),
			out2               => s_out2(7,23),
			lock_lower_row_out => s_locks_lower_out(7,23),
			lock_lower_row_in  => s_locks_lower_in(7,23),
			in1                => s_in1(7,23),
			in2                => s_in2(7,23),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(23)
		);
	s_in1(7,23)            <= s_out1(8,23);
	s_in2(7,23)            <= s_out2(8,24);
	s_locks_lower_in(7,23) <= s_locks_lower_out(8,23);

		normal_cell_7_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,24),
			fetch              => s_fetch(7,24),
			data_in            => s_data_in(7,24),
			data_out           => s_data_out(7,24),
			out1               => s_out1(7,24),
			out2               => s_out2(7,24),
			lock_lower_row_out => s_locks_lower_out(7,24),
			lock_lower_row_in  => s_locks_lower_in(7,24),
			in1                => s_in1(7,24),
			in2                => s_in2(7,24),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(24)
		);
	s_in1(7,24)            <= s_out1(8,24);
	s_in2(7,24)            <= s_out2(8,25);
	s_locks_lower_in(7,24) <= s_locks_lower_out(8,24);

		normal_cell_7_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,25),
			fetch              => s_fetch(7,25),
			data_in            => s_data_in(7,25),
			data_out           => s_data_out(7,25),
			out1               => s_out1(7,25),
			out2               => s_out2(7,25),
			lock_lower_row_out => s_locks_lower_out(7,25),
			lock_lower_row_in  => s_locks_lower_in(7,25),
			in1                => s_in1(7,25),
			in2                => s_in2(7,25),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(25)
		);
	s_in1(7,25)            <= s_out1(8,25);
	s_in2(7,25)            <= s_out2(8,26);
	s_locks_lower_in(7,25) <= s_locks_lower_out(8,25);

		normal_cell_7_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,26),
			fetch              => s_fetch(7,26),
			data_in            => s_data_in(7,26),
			data_out           => s_data_out(7,26),
			out1               => s_out1(7,26),
			out2               => s_out2(7,26),
			lock_lower_row_out => s_locks_lower_out(7,26),
			lock_lower_row_in  => s_locks_lower_in(7,26),
			in1                => s_in1(7,26),
			in2                => s_in2(7,26),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(26)
		);
	s_in1(7,26)            <= s_out1(8,26);
	s_in2(7,26)            <= s_out2(8,27);
	s_locks_lower_in(7,26) <= s_locks_lower_out(8,26);

		normal_cell_7_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,27),
			fetch              => s_fetch(7,27),
			data_in            => s_data_in(7,27),
			data_out           => s_data_out(7,27),
			out1               => s_out1(7,27),
			out2               => s_out2(7,27),
			lock_lower_row_out => s_locks_lower_out(7,27),
			lock_lower_row_in  => s_locks_lower_in(7,27),
			in1                => s_in1(7,27),
			in2                => s_in2(7,27),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(27)
		);
	s_in1(7,27)            <= s_out1(8,27);
	s_in2(7,27)            <= s_out2(8,28);
	s_locks_lower_in(7,27) <= s_locks_lower_out(8,27);

		normal_cell_7_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,28),
			fetch              => s_fetch(7,28),
			data_in            => s_data_in(7,28),
			data_out           => s_data_out(7,28),
			out1               => s_out1(7,28),
			out2               => s_out2(7,28),
			lock_lower_row_out => s_locks_lower_out(7,28),
			lock_lower_row_in  => s_locks_lower_in(7,28),
			in1                => s_in1(7,28),
			in2                => s_in2(7,28),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(28)
		);
	s_in1(7,28)            <= s_out1(8,28);
	s_in2(7,28)            <= s_out2(8,29);
	s_locks_lower_in(7,28) <= s_locks_lower_out(8,28);

		normal_cell_7_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,29),
			fetch              => s_fetch(7,29),
			data_in            => s_data_in(7,29),
			data_out           => s_data_out(7,29),
			out1               => s_out1(7,29),
			out2               => s_out2(7,29),
			lock_lower_row_out => s_locks_lower_out(7,29),
			lock_lower_row_in  => s_locks_lower_in(7,29),
			in1                => s_in1(7,29),
			in2                => s_in2(7,29),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(29)
		);
	s_in1(7,29)            <= s_out1(8,29);
	s_in2(7,29)            <= s_out2(8,30);
	s_locks_lower_in(7,29) <= s_locks_lower_out(8,29);

		normal_cell_7_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,30),
			fetch              => s_fetch(7,30),
			data_in            => s_data_in(7,30),
			data_out           => s_data_out(7,30),
			out1               => s_out1(7,30),
			out2               => s_out2(7,30),
			lock_lower_row_out => s_locks_lower_out(7,30),
			lock_lower_row_in  => s_locks_lower_in(7,30),
			in1                => s_in1(7,30),
			in2                => s_in2(7,30),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(30)
		);
	s_in1(7,30)            <= s_out1(8,30);
	s_in2(7,30)            <= s_out2(8,31);
	s_locks_lower_in(7,30) <= s_locks_lower_out(8,30);

		normal_cell_7_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,31),
			fetch              => s_fetch(7,31),
			data_in            => s_data_in(7,31),
			data_out           => s_data_out(7,31),
			out1               => s_out1(7,31),
			out2               => s_out2(7,31),
			lock_lower_row_out => s_locks_lower_out(7,31),
			lock_lower_row_in  => s_locks_lower_in(7,31),
			in1                => s_in1(7,31),
			in2                => s_in2(7,31),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(31)
		);
	s_in1(7,31)            <= s_out1(8,31);
	s_in2(7,31)            <= s_out2(8,32);
	s_locks_lower_in(7,31) <= s_locks_lower_out(8,31);

		normal_cell_7_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,32),
			fetch              => s_fetch(7,32),
			data_in            => s_data_in(7,32),
			data_out           => s_data_out(7,32),
			out1               => s_out1(7,32),
			out2               => s_out2(7,32),
			lock_lower_row_out => s_locks_lower_out(7,32),
			lock_lower_row_in  => s_locks_lower_in(7,32),
			in1                => s_in1(7,32),
			in2                => s_in2(7,32),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(32)
		);
	s_in1(7,32)            <= s_out1(8,32);
	s_in2(7,32)            <= s_out2(8,33);
	s_locks_lower_in(7,32) <= s_locks_lower_out(8,32);

		normal_cell_7_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,33),
			fetch              => s_fetch(7,33),
			data_in            => s_data_in(7,33),
			data_out           => s_data_out(7,33),
			out1               => s_out1(7,33),
			out2               => s_out2(7,33),
			lock_lower_row_out => s_locks_lower_out(7,33),
			lock_lower_row_in  => s_locks_lower_in(7,33),
			in1                => s_in1(7,33),
			in2                => s_in2(7,33),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(33)
		);
	s_in1(7,33)            <= s_out1(8,33);
	s_in2(7,33)            <= s_out2(8,34);
	s_locks_lower_in(7,33) <= s_locks_lower_out(8,33);

		normal_cell_7_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,34),
			fetch              => s_fetch(7,34),
			data_in            => s_data_in(7,34),
			data_out           => s_data_out(7,34),
			out1               => s_out1(7,34),
			out2               => s_out2(7,34),
			lock_lower_row_out => s_locks_lower_out(7,34),
			lock_lower_row_in  => s_locks_lower_in(7,34),
			in1                => s_in1(7,34),
			in2                => s_in2(7,34),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(34)
		);
	s_in1(7,34)            <= s_out1(8,34);
	s_in2(7,34)            <= s_out2(8,35);
	s_locks_lower_in(7,34) <= s_locks_lower_out(8,34);

		normal_cell_7_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,35),
			fetch              => s_fetch(7,35),
			data_in            => s_data_in(7,35),
			data_out           => s_data_out(7,35),
			out1               => s_out1(7,35),
			out2               => s_out2(7,35),
			lock_lower_row_out => s_locks_lower_out(7,35),
			lock_lower_row_in  => s_locks_lower_in(7,35),
			in1                => s_in1(7,35),
			in2                => s_in2(7,35),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(35)
		);
	s_in1(7,35)            <= s_out1(8,35);
	s_in2(7,35)            <= s_out2(8,36);
	s_locks_lower_in(7,35) <= s_locks_lower_out(8,35);

		normal_cell_7_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,36),
			fetch              => s_fetch(7,36),
			data_in            => s_data_in(7,36),
			data_out           => s_data_out(7,36),
			out1               => s_out1(7,36),
			out2               => s_out2(7,36),
			lock_lower_row_out => s_locks_lower_out(7,36),
			lock_lower_row_in  => s_locks_lower_in(7,36),
			in1                => s_in1(7,36),
			in2                => s_in2(7,36),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(36)
		);
	s_in1(7,36)            <= s_out1(8,36);
	s_in2(7,36)            <= s_out2(8,37);
	s_locks_lower_in(7,36) <= s_locks_lower_out(8,36);

		normal_cell_7_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,37),
			fetch              => s_fetch(7,37),
			data_in            => s_data_in(7,37),
			data_out           => s_data_out(7,37),
			out1               => s_out1(7,37),
			out2               => s_out2(7,37),
			lock_lower_row_out => s_locks_lower_out(7,37),
			lock_lower_row_in  => s_locks_lower_in(7,37),
			in1                => s_in1(7,37),
			in2                => s_in2(7,37),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(37)
		);
	s_in1(7,37)            <= s_out1(8,37);
	s_in2(7,37)            <= s_out2(8,38);
	s_locks_lower_in(7,37) <= s_locks_lower_out(8,37);

		normal_cell_7_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,38),
			fetch              => s_fetch(7,38),
			data_in            => s_data_in(7,38),
			data_out           => s_data_out(7,38),
			out1               => s_out1(7,38),
			out2               => s_out2(7,38),
			lock_lower_row_out => s_locks_lower_out(7,38),
			lock_lower_row_in  => s_locks_lower_in(7,38),
			in1                => s_in1(7,38),
			in2                => s_in2(7,38),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(38)
		);
	s_in1(7,38)            <= s_out1(8,38);
	s_in2(7,38)            <= s_out2(8,39);
	s_locks_lower_in(7,38) <= s_locks_lower_out(8,38);

		normal_cell_7_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,39),
			fetch              => s_fetch(7,39),
			data_in            => s_data_in(7,39),
			data_out           => s_data_out(7,39),
			out1               => s_out1(7,39),
			out2               => s_out2(7,39),
			lock_lower_row_out => s_locks_lower_out(7,39),
			lock_lower_row_in  => s_locks_lower_in(7,39),
			in1                => s_in1(7,39),
			in2                => s_in2(7,39),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(39)
		);
	s_in1(7,39)            <= s_out1(8,39);
	s_in2(7,39)            <= s_out2(8,40);
	s_locks_lower_in(7,39) <= s_locks_lower_out(8,39);

		normal_cell_7_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,40),
			fetch              => s_fetch(7,40),
			data_in            => s_data_in(7,40),
			data_out           => s_data_out(7,40),
			out1               => s_out1(7,40),
			out2               => s_out2(7,40),
			lock_lower_row_out => s_locks_lower_out(7,40),
			lock_lower_row_in  => s_locks_lower_in(7,40),
			in1                => s_in1(7,40),
			in2                => s_in2(7,40),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(40)
		);
	s_in1(7,40)            <= s_out1(8,40);
	s_in2(7,40)            <= s_out2(8,41);
	s_locks_lower_in(7,40) <= s_locks_lower_out(8,40);

		normal_cell_7_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,41),
			fetch              => s_fetch(7,41),
			data_in            => s_data_in(7,41),
			data_out           => s_data_out(7,41),
			out1               => s_out1(7,41),
			out2               => s_out2(7,41),
			lock_lower_row_out => s_locks_lower_out(7,41),
			lock_lower_row_in  => s_locks_lower_in(7,41),
			in1                => s_in1(7,41),
			in2                => s_in2(7,41),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(41)
		);
	s_in1(7,41)            <= s_out1(8,41);
	s_in2(7,41)            <= s_out2(8,42);
	s_locks_lower_in(7,41) <= s_locks_lower_out(8,41);

		normal_cell_7_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,42),
			fetch              => s_fetch(7,42),
			data_in            => s_data_in(7,42),
			data_out           => s_data_out(7,42),
			out1               => s_out1(7,42),
			out2               => s_out2(7,42),
			lock_lower_row_out => s_locks_lower_out(7,42),
			lock_lower_row_in  => s_locks_lower_in(7,42),
			in1                => s_in1(7,42),
			in2                => s_in2(7,42),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(42)
		);
	s_in1(7,42)            <= s_out1(8,42);
	s_in2(7,42)            <= s_out2(8,43);
	s_locks_lower_in(7,42) <= s_locks_lower_out(8,42);

		normal_cell_7_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,43),
			fetch              => s_fetch(7,43),
			data_in            => s_data_in(7,43),
			data_out           => s_data_out(7,43),
			out1               => s_out1(7,43),
			out2               => s_out2(7,43),
			lock_lower_row_out => s_locks_lower_out(7,43),
			lock_lower_row_in  => s_locks_lower_in(7,43),
			in1                => s_in1(7,43),
			in2                => s_in2(7,43),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(43)
		);
	s_in1(7,43)            <= s_out1(8,43);
	s_in2(7,43)            <= s_out2(8,44);
	s_locks_lower_in(7,43) <= s_locks_lower_out(8,43);

		normal_cell_7_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,44),
			fetch              => s_fetch(7,44),
			data_in            => s_data_in(7,44),
			data_out           => s_data_out(7,44),
			out1               => s_out1(7,44),
			out2               => s_out2(7,44),
			lock_lower_row_out => s_locks_lower_out(7,44),
			lock_lower_row_in  => s_locks_lower_in(7,44),
			in1                => s_in1(7,44),
			in2                => s_in2(7,44),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(44)
		);
	s_in1(7,44)            <= s_out1(8,44);
	s_in2(7,44)            <= s_out2(8,45);
	s_locks_lower_in(7,44) <= s_locks_lower_out(8,44);

		normal_cell_7_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,45),
			fetch              => s_fetch(7,45),
			data_in            => s_data_in(7,45),
			data_out           => s_data_out(7,45),
			out1               => s_out1(7,45),
			out2               => s_out2(7,45),
			lock_lower_row_out => s_locks_lower_out(7,45),
			lock_lower_row_in  => s_locks_lower_in(7,45),
			in1                => s_in1(7,45),
			in2                => s_in2(7,45),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(45)
		);
	s_in1(7,45)            <= s_out1(8,45);
	s_in2(7,45)            <= s_out2(8,46);
	s_locks_lower_in(7,45) <= s_locks_lower_out(8,45);

		normal_cell_7_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,46),
			fetch              => s_fetch(7,46),
			data_in            => s_data_in(7,46),
			data_out           => s_data_out(7,46),
			out1               => s_out1(7,46),
			out2               => s_out2(7,46),
			lock_lower_row_out => s_locks_lower_out(7,46),
			lock_lower_row_in  => s_locks_lower_in(7,46),
			in1                => s_in1(7,46),
			in2                => s_in2(7,46),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(46)
		);
	s_in1(7,46)            <= s_out1(8,46);
	s_in2(7,46)            <= s_out2(8,47);
	s_locks_lower_in(7,46) <= s_locks_lower_out(8,46);

		normal_cell_7_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,47),
			fetch              => s_fetch(7,47),
			data_in            => s_data_in(7,47),
			data_out           => s_data_out(7,47),
			out1               => s_out1(7,47),
			out2               => s_out2(7,47),
			lock_lower_row_out => s_locks_lower_out(7,47),
			lock_lower_row_in  => s_locks_lower_in(7,47),
			in1                => s_in1(7,47),
			in2                => s_in2(7,47),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(47)
		);
	s_in1(7,47)            <= s_out1(8,47);
	s_in2(7,47)            <= s_out2(8,48);
	s_locks_lower_in(7,47) <= s_locks_lower_out(8,47);

		normal_cell_7_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,48),
			fetch              => s_fetch(7,48),
			data_in            => s_data_in(7,48),
			data_out           => s_data_out(7,48),
			out1               => s_out1(7,48),
			out2               => s_out2(7,48),
			lock_lower_row_out => s_locks_lower_out(7,48),
			lock_lower_row_in  => s_locks_lower_in(7,48),
			in1                => s_in1(7,48),
			in2                => s_in2(7,48),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(48)
		);
	s_in1(7,48)            <= s_out1(8,48);
	s_in2(7,48)            <= s_out2(8,49);
	s_locks_lower_in(7,48) <= s_locks_lower_out(8,48);

		normal_cell_7_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,49),
			fetch              => s_fetch(7,49),
			data_in            => s_data_in(7,49),
			data_out           => s_data_out(7,49),
			out1               => s_out1(7,49),
			out2               => s_out2(7,49),
			lock_lower_row_out => s_locks_lower_out(7,49),
			lock_lower_row_in  => s_locks_lower_in(7,49),
			in1                => s_in1(7,49),
			in2                => s_in2(7,49),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(49)
		);
	s_in1(7,49)            <= s_out1(8,49);
	s_in2(7,49)            <= s_out2(8,50);
	s_locks_lower_in(7,49) <= s_locks_lower_out(8,49);

		normal_cell_7_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,50),
			fetch              => s_fetch(7,50),
			data_in            => s_data_in(7,50),
			data_out           => s_data_out(7,50),
			out1               => s_out1(7,50),
			out2               => s_out2(7,50),
			lock_lower_row_out => s_locks_lower_out(7,50),
			lock_lower_row_in  => s_locks_lower_in(7,50),
			in1                => s_in1(7,50),
			in2                => s_in2(7,50),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(50)
		);
	s_in1(7,50)            <= s_out1(8,50);
	s_in2(7,50)            <= s_out2(8,51);
	s_locks_lower_in(7,50) <= s_locks_lower_out(8,50);

		normal_cell_7_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,51),
			fetch              => s_fetch(7,51),
			data_in            => s_data_in(7,51),
			data_out           => s_data_out(7,51),
			out1               => s_out1(7,51),
			out2               => s_out2(7,51),
			lock_lower_row_out => s_locks_lower_out(7,51),
			lock_lower_row_in  => s_locks_lower_in(7,51),
			in1                => s_in1(7,51),
			in2                => s_in2(7,51),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(51)
		);
	s_in1(7,51)            <= s_out1(8,51);
	s_in2(7,51)            <= s_out2(8,52);
	s_locks_lower_in(7,51) <= s_locks_lower_out(8,51);

		normal_cell_7_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,52),
			fetch              => s_fetch(7,52),
			data_in            => s_data_in(7,52),
			data_out           => s_data_out(7,52),
			out1               => s_out1(7,52),
			out2               => s_out2(7,52),
			lock_lower_row_out => s_locks_lower_out(7,52),
			lock_lower_row_in  => s_locks_lower_in(7,52),
			in1                => s_in1(7,52),
			in2                => s_in2(7,52),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(52)
		);
	s_in1(7,52)            <= s_out1(8,52);
	s_in2(7,52)            <= s_out2(8,53);
	s_locks_lower_in(7,52) <= s_locks_lower_out(8,52);

		normal_cell_7_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,53),
			fetch              => s_fetch(7,53),
			data_in            => s_data_in(7,53),
			data_out           => s_data_out(7,53),
			out1               => s_out1(7,53),
			out2               => s_out2(7,53),
			lock_lower_row_out => s_locks_lower_out(7,53),
			lock_lower_row_in  => s_locks_lower_in(7,53),
			in1                => s_in1(7,53),
			in2                => s_in2(7,53),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(53)
		);
	s_in1(7,53)            <= s_out1(8,53);
	s_in2(7,53)            <= s_out2(8,54);
	s_locks_lower_in(7,53) <= s_locks_lower_out(8,53);

		normal_cell_7_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,54),
			fetch              => s_fetch(7,54),
			data_in            => s_data_in(7,54),
			data_out           => s_data_out(7,54),
			out1               => s_out1(7,54),
			out2               => s_out2(7,54),
			lock_lower_row_out => s_locks_lower_out(7,54),
			lock_lower_row_in  => s_locks_lower_in(7,54),
			in1                => s_in1(7,54),
			in2                => s_in2(7,54),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(54)
		);
	s_in1(7,54)            <= s_out1(8,54);
	s_in2(7,54)            <= s_out2(8,55);
	s_locks_lower_in(7,54) <= s_locks_lower_out(8,54);

		normal_cell_7_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,55),
			fetch              => s_fetch(7,55),
			data_in            => s_data_in(7,55),
			data_out           => s_data_out(7,55),
			out1               => s_out1(7,55),
			out2               => s_out2(7,55),
			lock_lower_row_out => s_locks_lower_out(7,55),
			lock_lower_row_in  => s_locks_lower_in(7,55),
			in1                => s_in1(7,55),
			in2                => s_in2(7,55),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(55)
		);
	s_in1(7,55)            <= s_out1(8,55);
	s_in2(7,55)            <= s_out2(8,56);
	s_locks_lower_in(7,55) <= s_locks_lower_out(8,55);

		normal_cell_7_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,56),
			fetch              => s_fetch(7,56),
			data_in            => s_data_in(7,56),
			data_out           => s_data_out(7,56),
			out1               => s_out1(7,56),
			out2               => s_out2(7,56),
			lock_lower_row_out => s_locks_lower_out(7,56),
			lock_lower_row_in  => s_locks_lower_in(7,56),
			in1                => s_in1(7,56),
			in2                => s_in2(7,56),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(56)
		);
	s_in1(7,56)            <= s_out1(8,56);
	s_in2(7,56)            <= s_out2(8,57);
	s_locks_lower_in(7,56) <= s_locks_lower_out(8,56);

		normal_cell_7_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,57),
			fetch              => s_fetch(7,57),
			data_in            => s_data_in(7,57),
			data_out           => s_data_out(7,57),
			out1               => s_out1(7,57),
			out2               => s_out2(7,57),
			lock_lower_row_out => s_locks_lower_out(7,57),
			lock_lower_row_in  => s_locks_lower_in(7,57),
			in1                => s_in1(7,57),
			in2                => s_in2(7,57),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(57)
		);
	s_in1(7,57)            <= s_out1(8,57);
	s_in2(7,57)            <= s_out2(8,58);
	s_locks_lower_in(7,57) <= s_locks_lower_out(8,57);

		normal_cell_7_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,58),
			fetch              => s_fetch(7,58),
			data_in            => s_data_in(7,58),
			data_out           => s_data_out(7,58),
			out1               => s_out1(7,58),
			out2               => s_out2(7,58),
			lock_lower_row_out => s_locks_lower_out(7,58),
			lock_lower_row_in  => s_locks_lower_in(7,58),
			in1                => s_in1(7,58),
			in2                => s_in2(7,58),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(58)
		);
	s_in1(7,58)            <= s_out1(8,58);
	s_in2(7,58)            <= s_out2(8,59);
	s_locks_lower_in(7,58) <= s_locks_lower_out(8,58);

		normal_cell_7_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,59),
			fetch              => s_fetch(7,59),
			data_in            => s_data_in(7,59),
			data_out           => s_data_out(7,59),
			out1               => s_out1(7,59),
			out2               => s_out2(7,59),
			lock_lower_row_out => s_locks_lower_out(7,59),
			lock_lower_row_in  => s_locks_lower_in(7,59),
			in1                => s_in1(7,59),
			in2                => s_in2(7,59),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(59)
		);
	s_in1(7,59)            <= s_out1(8,59);
	s_in2(7,59)            <= s_out2(8,60);
	s_locks_lower_in(7,59) <= s_locks_lower_out(8,59);

		last_col_cell_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(7,60),
			fetch              => s_fetch(7,60),
			data_in            => s_data_in(7,60),
			data_out           => s_data_out(7,60),
			out1               => s_out1(7,60),
			out2               => s_out2(7,60),
			lock_lower_row_out => s_locks_lower_out(7,60),
			lock_lower_row_in  => s_locks_lower_in(7,60),
			in1                => s_in1(7,60),
			in2                => (others => '0'),
			lock_row           => s_locks(7),
			piv_found          => s_piv_found,
			row_data           => s_row_data(7),
			col_data           => s_col_data(60)
		);
	s_in1(7,60)            <= s_out1(8,60);
	s_locks_lower_in(7,60) <= s_locks_lower_out(8,60);

		normal_cell_8_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,1),
			fetch              => s_fetch(8,1),
			data_in            => s_data_in(8,1),
			data_out           => s_data_out(8,1),
			out1               => s_out1(8,1),
			out2               => s_out2(8,1),
			lock_lower_row_out => s_locks_lower_out(8,1),
			lock_lower_row_in  => s_locks_lower_in(8,1),
			in1                => s_in1(8,1),
			in2                => s_in2(8,1),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(1)
		);
	s_in1(8,1)            <= s_out1(9,1);
	s_in2(8,1)            <= s_out2(9,2);
	s_locks_lower_in(8,1) <= s_locks_lower_out(9,1);

		normal_cell_8_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,2),
			fetch              => s_fetch(8,2),
			data_in            => s_data_in(8,2),
			data_out           => s_data_out(8,2),
			out1               => s_out1(8,2),
			out2               => s_out2(8,2),
			lock_lower_row_out => s_locks_lower_out(8,2),
			lock_lower_row_in  => s_locks_lower_in(8,2),
			in1                => s_in1(8,2),
			in2                => s_in2(8,2),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(2)
		);
	s_in1(8,2)            <= s_out1(9,2);
	s_in2(8,2)            <= s_out2(9,3);
	s_locks_lower_in(8,2) <= s_locks_lower_out(9,2);

		normal_cell_8_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,3),
			fetch              => s_fetch(8,3),
			data_in            => s_data_in(8,3),
			data_out           => s_data_out(8,3),
			out1               => s_out1(8,3),
			out2               => s_out2(8,3),
			lock_lower_row_out => s_locks_lower_out(8,3),
			lock_lower_row_in  => s_locks_lower_in(8,3),
			in1                => s_in1(8,3),
			in2                => s_in2(8,3),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(3)
		);
	s_in1(8,3)            <= s_out1(9,3);
	s_in2(8,3)            <= s_out2(9,4);
	s_locks_lower_in(8,3) <= s_locks_lower_out(9,3);

		normal_cell_8_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,4),
			fetch              => s_fetch(8,4),
			data_in            => s_data_in(8,4),
			data_out           => s_data_out(8,4),
			out1               => s_out1(8,4),
			out2               => s_out2(8,4),
			lock_lower_row_out => s_locks_lower_out(8,4),
			lock_lower_row_in  => s_locks_lower_in(8,4),
			in1                => s_in1(8,4),
			in2                => s_in2(8,4),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(4)
		);
	s_in1(8,4)            <= s_out1(9,4);
	s_in2(8,4)            <= s_out2(9,5);
	s_locks_lower_in(8,4) <= s_locks_lower_out(9,4);

		normal_cell_8_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,5),
			fetch              => s_fetch(8,5),
			data_in            => s_data_in(8,5),
			data_out           => s_data_out(8,5),
			out1               => s_out1(8,5),
			out2               => s_out2(8,5),
			lock_lower_row_out => s_locks_lower_out(8,5),
			lock_lower_row_in  => s_locks_lower_in(8,5),
			in1                => s_in1(8,5),
			in2                => s_in2(8,5),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(5)
		);
	s_in1(8,5)            <= s_out1(9,5);
	s_in2(8,5)            <= s_out2(9,6);
	s_locks_lower_in(8,5) <= s_locks_lower_out(9,5);

		normal_cell_8_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,6),
			fetch              => s_fetch(8,6),
			data_in            => s_data_in(8,6),
			data_out           => s_data_out(8,6),
			out1               => s_out1(8,6),
			out2               => s_out2(8,6),
			lock_lower_row_out => s_locks_lower_out(8,6),
			lock_lower_row_in  => s_locks_lower_in(8,6),
			in1                => s_in1(8,6),
			in2                => s_in2(8,6),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(6)
		);
	s_in1(8,6)            <= s_out1(9,6);
	s_in2(8,6)            <= s_out2(9,7);
	s_locks_lower_in(8,6) <= s_locks_lower_out(9,6);

		normal_cell_8_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,7),
			fetch              => s_fetch(8,7),
			data_in            => s_data_in(8,7),
			data_out           => s_data_out(8,7),
			out1               => s_out1(8,7),
			out2               => s_out2(8,7),
			lock_lower_row_out => s_locks_lower_out(8,7),
			lock_lower_row_in  => s_locks_lower_in(8,7),
			in1                => s_in1(8,7),
			in2                => s_in2(8,7),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(7)
		);
	s_in1(8,7)            <= s_out1(9,7);
	s_in2(8,7)            <= s_out2(9,8);
	s_locks_lower_in(8,7) <= s_locks_lower_out(9,7);

		normal_cell_8_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,8),
			fetch              => s_fetch(8,8),
			data_in            => s_data_in(8,8),
			data_out           => s_data_out(8,8),
			out1               => s_out1(8,8),
			out2               => s_out2(8,8),
			lock_lower_row_out => s_locks_lower_out(8,8),
			lock_lower_row_in  => s_locks_lower_in(8,8),
			in1                => s_in1(8,8),
			in2                => s_in2(8,8),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(8)
		);
	s_in1(8,8)            <= s_out1(9,8);
	s_in2(8,8)            <= s_out2(9,9);
	s_locks_lower_in(8,8) <= s_locks_lower_out(9,8);

		normal_cell_8_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,9),
			fetch              => s_fetch(8,9),
			data_in            => s_data_in(8,9),
			data_out           => s_data_out(8,9),
			out1               => s_out1(8,9),
			out2               => s_out2(8,9),
			lock_lower_row_out => s_locks_lower_out(8,9),
			lock_lower_row_in  => s_locks_lower_in(8,9),
			in1                => s_in1(8,9),
			in2                => s_in2(8,9),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(9)
		);
	s_in1(8,9)            <= s_out1(9,9);
	s_in2(8,9)            <= s_out2(9,10);
	s_locks_lower_in(8,9) <= s_locks_lower_out(9,9);

		normal_cell_8_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,10),
			fetch              => s_fetch(8,10),
			data_in            => s_data_in(8,10),
			data_out           => s_data_out(8,10),
			out1               => s_out1(8,10),
			out2               => s_out2(8,10),
			lock_lower_row_out => s_locks_lower_out(8,10),
			lock_lower_row_in  => s_locks_lower_in(8,10),
			in1                => s_in1(8,10),
			in2                => s_in2(8,10),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(10)
		);
	s_in1(8,10)            <= s_out1(9,10);
	s_in2(8,10)            <= s_out2(9,11);
	s_locks_lower_in(8,10) <= s_locks_lower_out(9,10);

		normal_cell_8_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,11),
			fetch              => s_fetch(8,11),
			data_in            => s_data_in(8,11),
			data_out           => s_data_out(8,11),
			out1               => s_out1(8,11),
			out2               => s_out2(8,11),
			lock_lower_row_out => s_locks_lower_out(8,11),
			lock_lower_row_in  => s_locks_lower_in(8,11),
			in1                => s_in1(8,11),
			in2                => s_in2(8,11),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(11)
		);
	s_in1(8,11)            <= s_out1(9,11);
	s_in2(8,11)            <= s_out2(9,12);
	s_locks_lower_in(8,11) <= s_locks_lower_out(9,11);

		normal_cell_8_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,12),
			fetch              => s_fetch(8,12),
			data_in            => s_data_in(8,12),
			data_out           => s_data_out(8,12),
			out1               => s_out1(8,12),
			out2               => s_out2(8,12),
			lock_lower_row_out => s_locks_lower_out(8,12),
			lock_lower_row_in  => s_locks_lower_in(8,12),
			in1                => s_in1(8,12),
			in2                => s_in2(8,12),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(12)
		);
	s_in1(8,12)            <= s_out1(9,12);
	s_in2(8,12)            <= s_out2(9,13);
	s_locks_lower_in(8,12) <= s_locks_lower_out(9,12);

		normal_cell_8_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,13),
			fetch              => s_fetch(8,13),
			data_in            => s_data_in(8,13),
			data_out           => s_data_out(8,13),
			out1               => s_out1(8,13),
			out2               => s_out2(8,13),
			lock_lower_row_out => s_locks_lower_out(8,13),
			lock_lower_row_in  => s_locks_lower_in(8,13),
			in1                => s_in1(8,13),
			in2                => s_in2(8,13),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(13)
		);
	s_in1(8,13)            <= s_out1(9,13);
	s_in2(8,13)            <= s_out2(9,14);
	s_locks_lower_in(8,13) <= s_locks_lower_out(9,13);

		normal_cell_8_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,14),
			fetch              => s_fetch(8,14),
			data_in            => s_data_in(8,14),
			data_out           => s_data_out(8,14),
			out1               => s_out1(8,14),
			out2               => s_out2(8,14),
			lock_lower_row_out => s_locks_lower_out(8,14),
			lock_lower_row_in  => s_locks_lower_in(8,14),
			in1                => s_in1(8,14),
			in2                => s_in2(8,14),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(14)
		);
	s_in1(8,14)            <= s_out1(9,14);
	s_in2(8,14)            <= s_out2(9,15);
	s_locks_lower_in(8,14) <= s_locks_lower_out(9,14);

		normal_cell_8_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,15),
			fetch              => s_fetch(8,15),
			data_in            => s_data_in(8,15),
			data_out           => s_data_out(8,15),
			out1               => s_out1(8,15),
			out2               => s_out2(8,15),
			lock_lower_row_out => s_locks_lower_out(8,15),
			lock_lower_row_in  => s_locks_lower_in(8,15),
			in1                => s_in1(8,15),
			in2                => s_in2(8,15),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(15)
		);
	s_in1(8,15)            <= s_out1(9,15);
	s_in2(8,15)            <= s_out2(9,16);
	s_locks_lower_in(8,15) <= s_locks_lower_out(9,15);

		normal_cell_8_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,16),
			fetch              => s_fetch(8,16),
			data_in            => s_data_in(8,16),
			data_out           => s_data_out(8,16),
			out1               => s_out1(8,16),
			out2               => s_out2(8,16),
			lock_lower_row_out => s_locks_lower_out(8,16),
			lock_lower_row_in  => s_locks_lower_in(8,16),
			in1                => s_in1(8,16),
			in2                => s_in2(8,16),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(16)
		);
	s_in1(8,16)            <= s_out1(9,16);
	s_in2(8,16)            <= s_out2(9,17);
	s_locks_lower_in(8,16) <= s_locks_lower_out(9,16);

		normal_cell_8_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,17),
			fetch              => s_fetch(8,17),
			data_in            => s_data_in(8,17),
			data_out           => s_data_out(8,17),
			out1               => s_out1(8,17),
			out2               => s_out2(8,17),
			lock_lower_row_out => s_locks_lower_out(8,17),
			lock_lower_row_in  => s_locks_lower_in(8,17),
			in1                => s_in1(8,17),
			in2                => s_in2(8,17),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(17)
		);
	s_in1(8,17)            <= s_out1(9,17);
	s_in2(8,17)            <= s_out2(9,18);
	s_locks_lower_in(8,17) <= s_locks_lower_out(9,17);

		normal_cell_8_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,18),
			fetch              => s_fetch(8,18),
			data_in            => s_data_in(8,18),
			data_out           => s_data_out(8,18),
			out1               => s_out1(8,18),
			out2               => s_out2(8,18),
			lock_lower_row_out => s_locks_lower_out(8,18),
			lock_lower_row_in  => s_locks_lower_in(8,18),
			in1                => s_in1(8,18),
			in2                => s_in2(8,18),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(18)
		);
	s_in1(8,18)            <= s_out1(9,18);
	s_in2(8,18)            <= s_out2(9,19);
	s_locks_lower_in(8,18) <= s_locks_lower_out(9,18);

		normal_cell_8_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,19),
			fetch              => s_fetch(8,19),
			data_in            => s_data_in(8,19),
			data_out           => s_data_out(8,19),
			out1               => s_out1(8,19),
			out2               => s_out2(8,19),
			lock_lower_row_out => s_locks_lower_out(8,19),
			lock_lower_row_in  => s_locks_lower_in(8,19),
			in1                => s_in1(8,19),
			in2                => s_in2(8,19),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(19)
		);
	s_in1(8,19)            <= s_out1(9,19);
	s_in2(8,19)            <= s_out2(9,20);
	s_locks_lower_in(8,19) <= s_locks_lower_out(9,19);

		normal_cell_8_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,20),
			fetch              => s_fetch(8,20),
			data_in            => s_data_in(8,20),
			data_out           => s_data_out(8,20),
			out1               => s_out1(8,20),
			out2               => s_out2(8,20),
			lock_lower_row_out => s_locks_lower_out(8,20),
			lock_lower_row_in  => s_locks_lower_in(8,20),
			in1                => s_in1(8,20),
			in2                => s_in2(8,20),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(20)
		);
	s_in1(8,20)            <= s_out1(9,20);
	s_in2(8,20)            <= s_out2(9,21);
	s_locks_lower_in(8,20) <= s_locks_lower_out(9,20);

		normal_cell_8_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,21),
			fetch              => s_fetch(8,21),
			data_in            => s_data_in(8,21),
			data_out           => s_data_out(8,21),
			out1               => s_out1(8,21),
			out2               => s_out2(8,21),
			lock_lower_row_out => s_locks_lower_out(8,21),
			lock_lower_row_in  => s_locks_lower_in(8,21),
			in1                => s_in1(8,21),
			in2                => s_in2(8,21),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(21)
		);
	s_in1(8,21)            <= s_out1(9,21);
	s_in2(8,21)            <= s_out2(9,22);
	s_locks_lower_in(8,21) <= s_locks_lower_out(9,21);

		normal_cell_8_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,22),
			fetch              => s_fetch(8,22),
			data_in            => s_data_in(8,22),
			data_out           => s_data_out(8,22),
			out1               => s_out1(8,22),
			out2               => s_out2(8,22),
			lock_lower_row_out => s_locks_lower_out(8,22),
			lock_lower_row_in  => s_locks_lower_in(8,22),
			in1                => s_in1(8,22),
			in2                => s_in2(8,22),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(22)
		);
	s_in1(8,22)            <= s_out1(9,22);
	s_in2(8,22)            <= s_out2(9,23);
	s_locks_lower_in(8,22) <= s_locks_lower_out(9,22);

		normal_cell_8_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,23),
			fetch              => s_fetch(8,23),
			data_in            => s_data_in(8,23),
			data_out           => s_data_out(8,23),
			out1               => s_out1(8,23),
			out2               => s_out2(8,23),
			lock_lower_row_out => s_locks_lower_out(8,23),
			lock_lower_row_in  => s_locks_lower_in(8,23),
			in1                => s_in1(8,23),
			in2                => s_in2(8,23),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(23)
		);
	s_in1(8,23)            <= s_out1(9,23);
	s_in2(8,23)            <= s_out2(9,24);
	s_locks_lower_in(8,23) <= s_locks_lower_out(9,23);

		normal_cell_8_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,24),
			fetch              => s_fetch(8,24),
			data_in            => s_data_in(8,24),
			data_out           => s_data_out(8,24),
			out1               => s_out1(8,24),
			out2               => s_out2(8,24),
			lock_lower_row_out => s_locks_lower_out(8,24),
			lock_lower_row_in  => s_locks_lower_in(8,24),
			in1                => s_in1(8,24),
			in2                => s_in2(8,24),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(24)
		);
	s_in1(8,24)            <= s_out1(9,24);
	s_in2(8,24)            <= s_out2(9,25);
	s_locks_lower_in(8,24) <= s_locks_lower_out(9,24);

		normal_cell_8_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,25),
			fetch              => s_fetch(8,25),
			data_in            => s_data_in(8,25),
			data_out           => s_data_out(8,25),
			out1               => s_out1(8,25),
			out2               => s_out2(8,25),
			lock_lower_row_out => s_locks_lower_out(8,25),
			lock_lower_row_in  => s_locks_lower_in(8,25),
			in1                => s_in1(8,25),
			in2                => s_in2(8,25),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(25)
		);
	s_in1(8,25)            <= s_out1(9,25);
	s_in2(8,25)            <= s_out2(9,26);
	s_locks_lower_in(8,25) <= s_locks_lower_out(9,25);

		normal_cell_8_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,26),
			fetch              => s_fetch(8,26),
			data_in            => s_data_in(8,26),
			data_out           => s_data_out(8,26),
			out1               => s_out1(8,26),
			out2               => s_out2(8,26),
			lock_lower_row_out => s_locks_lower_out(8,26),
			lock_lower_row_in  => s_locks_lower_in(8,26),
			in1                => s_in1(8,26),
			in2                => s_in2(8,26),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(26)
		);
	s_in1(8,26)            <= s_out1(9,26);
	s_in2(8,26)            <= s_out2(9,27);
	s_locks_lower_in(8,26) <= s_locks_lower_out(9,26);

		normal_cell_8_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,27),
			fetch              => s_fetch(8,27),
			data_in            => s_data_in(8,27),
			data_out           => s_data_out(8,27),
			out1               => s_out1(8,27),
			out2               => s_out2(8,27),
			lock_lower_row_out => s_locks_lower_out(8,27),
			lock_lower_row_in  => s_locks_lower_in(8,27),
			in1                => s_in1(8,27),
			in2                => s_in2(8,27),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(27)
		);
	s_in1(8,27)            <= s_out1(9,27);
	s_in2(8,27)            <= s_out2(9,28);
	s_locks_lower_in(8,27) <= s_locks_lower_out(9,27);

		normal_cell_8_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,28),
			fetch              => s_fetch(8,28),
			data_in            => s_data_in(8,28),
			data_out           => s_data_out(8,28),
			out1               => s_out1(8,28),
			out2               => s_out2(8,28),
			lock_lower_row_out => s_locks_lower_out(8,28),
			lock_lower_row_in  => s_locks_lower_in(8,28),
			in1                => s_in1(8,28),
			in2                => s_in2(8,28),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(28)
		);
	s_in1(8,28)            <= s_out1(9,28);
	s_in2(8,28)            <= s_out2(9,29);
	s_locks_lower_in(8,28) <= s_locks_lower_out(9,28);

		normal_cell_8_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,29),
			fetch              => s_fetch(8,29),
			data_in            => s_data_in(8,29),
			data_out           => s_data_out(8,29),
			out1               => s_out1(8,29),
			out2               => s_out2(8,29),
			lock_lower_row_out => s_locks_lower_out(8,29),
			lock_lower_row_in  => s_locks_lower_in(8,29),
			in1                => s_in1(8,29),
			in2                => s_in2(8,29),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(29)
		);
	s_in1(8,29)            <= s_out1(9,29);
	s_in2(8,29)            <= s_out2(9,30);
	s_locks_lower_in(8,29) <= s_locks_lower_out(9,29);

		normal_cell_8_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,30),
			fetch              => s_fetch(8,30),
			data_in            => s_data_in(8,30),
			data_out           => s_data_out(8,30),
			out1               => s_out1(8,30),
			out2               => s_out2(8,30),
			lock_lower_row_out => s_locks_lower_out(8,30),
			lock_lower_row_in  => s_locks_lower_in(8,30),
			in1                => s_in1(8,30),
			in2                => s_in2(8,30),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(30)
		);
	s_in1(8,30)            <= s_out1(9,30);
	s_in2(8,30)            <= s_out2(9,31);
	s_locks_lower_in(8,30) <= s_locks_lower_out(9,30);

		normal_cell_8_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,31),
			fetch              => s_fetch(8,31),
			data_in            => s_data_in(8,31),
			data_out           => s_data_out(8,31),
			out1               => s_out1(8,31),
			out2               => s_out2(8,31),
			lock_lower_row_out => s_locks_lower_out(8,31),
			lock_lower_row_in  => s_locks_lower_in(8,31),
			in1                => s_in1(8,31),
			in2                => s_in2(8,31),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(31)
		);
	s_in1(8,31)            <= s_out1(9,31);
	s_in2(8,31)            <= s_out2(9,32);
	s_locks_lower_in(8,31) <= s_locks_lower_out(9,31);

		normal_cell_8_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,32),
			fetch              => s_fetch(8,32),
			data_in            => s_data_in(8,32),
			data_out           => s_data_out(8,32),
			out1               => s_out1(8,32),
			out2               => s_out2(8,32),
			lock_lower_row_out => s_locks_lower_out(8,32),
			lock_lower_row_in  => s_locks_lower_in(8,32),
			in1                => s_in1(8,32),
			in2                => s_in2(8,32),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(32)
		);
	s_in1(8,32)            <= s_out1(9,32);
	s_in2(8,32)            <= s_out2(9,33);
	s_locks_lower_in(8,32) <= s_locks_lower_out(9,32);

		normal_cell_8_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,33),
			fetch              => s_fetch(8,33),
			data_in            => s_data_in(8,33),
			data_out           => s_data_out(8,33),
			out1               => s_out1(8,33),
			out2               => s_out2(8,33),
			lock_lower_row_out => s_locks_lower_out(8,33),
			lock_lower_row_in  => s_locks_lower_in(8,33),
			in1                => s_in1(8,33),
			in2                => s_in2(8,33),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(33)
		);
	s_in1(8,33)            <= s_out1(9,33);
	s_in2(8,33)            <= s_out2(9,34);
	s_locks_lower_in(8,33) <= s_locks_lower_out(9,33);

		normal_cell_8_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,34),
			fetch              => s_fetch(8,34),
			data_in            => s_data_in(8,34),
			data_out           => s_data_out(8,34),
			out1               => s_out1(8,34),
			out2               => s_out2(8,34),
			lock_lower_row_out => s_locks_lower_out(8,34),
			lock_lower_row_in  => s_locks_lower_in(8,34),
			in1                => s_in1(8,34),
			in2                => s_in2(8,34),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(34)
		);
	s_in1(8,34)            <= s_out1(9,34);
	s_in2(8,34)            <= s_out2(9,35);
	s_locks_lower_in(8,34) <= s_locks_lower_out(9,34);

		normal_cell_8_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,35),
			fetch              => s_fetch(8,35),
			data_in            => s_data_in(8,35),
			data_out           => s_data_out(8,35),
			out1               => s_out1(8,35),
			out2               => s_out2(8,35),
			lock_lower_row_out => s_locks_lower_out(8,35),
			lock_lower_row_in  => s_locks_lower_in(8,35),
			in1                => s_in1(8,35),
			in2                => s_in2(8,35),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(35)
		);
	s_in1(8,35)            <= s_out1(9,35);
	s_in2(8,35)            <= s_out2(9,36);
	s_locks_lower_in(8,35) <= s_locks_lower_out(9,35);

		normal_cell_8_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,36),
			fetch              => s_fetch(8,36),
			data_in            => s_data_in(8,36),
			data_out           => s_data_out(8,36),
			out1               => s_out1(8,36),
			out2               => s_out2(8,36),
			lock_lower_row_out => s_locks_lower_out(8,36),
			lock_lower_row_in  => s_locks_lower_in(8,36),
			in1                => s_in1(8,36),
			in2                => s_in2(8,36),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(36)
		);
	s_in1(8,36)            <= s_out1(9,36);
	s_in2(8,36)            <= s_out2(9,37);
	s_locks_lower_in(8,36) <= s_locks_lower_out(9,36);

		normal_cell_8_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,37),
			fetch              => s_fetch(8,37),
			data_in            => s_data_in(8,37),
			data_out           => s_data_out(8,37),
			out1               => s_out1(8,37),
			out2               => s_out2(8,37),
			lock_lower_row_out => s_locks_lower_out(8,37),
			lock_lower_row_in  => s_locks_lower_in(8,37),
			in1                => s_in1(8,37),
			in2                => s_in2(8,37),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(37)
		);
	s_in1(8,37)            <= s_out1(9,37);
	s_in2(8,37)            <= s_out2(9,38);
	s_locks_lower_in(8,37) <= s_locks_lower_out(9,37);

		normal_cell_8_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,38),
			fetch              => s_fetch(8,38),
			data_in            => s_data_in(8,38),
			data_out           => s_data_out(8,38),
			out1               => s_out1(8,38),
			out2               => s_out2(8,38),
			lock_lower_row_out => s_locks_lower_out(8,38),
			lock_lower_row_in  => s_locks_lower_in(8,38),
			in1                => s_in1(8,38),
			in2                => s_in2(8,38),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(38)
		);
	s_in1(8,38)            <= s_out1(9,38);
	s_in2(8,38)            <= s_out2(9,39);
	s_locks_lower_in(8,38) <= s_locks_lower_out(9,38);

		normal_cell_8_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,39),
			fetch              => s_fetch(8,39),
			data_in            => s_data_in(8,39),
			data_out           => s_data_out(8,39),
			out1               => s_out1(8,39),
			out2               => s_out2(8,39),
			lock_lower_row_out => s_locks_lower_out(8,39),
			lock_lower_row_in  => s_locks_lower_in(8,39),
			in1                => s_in1(8,39),
			in2                => s_in2(8,39),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(39)
		);
	s_in1(8,39)            <= s_out1(9,39);
	s_in2(8,39)            <= s_out2(9,40);
	s_locks_lower_in(8,39) <= s_locks_lower_out(9,39);

		normal_cell_8_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,40),
			fetch              => s_fetch(8,40),
			data_in            => s_data_in(8,40),
			data_out           => s_data_out(8,40),
			out1               => s_out1(8,40),
			out2               => s_out2(8,40),
			lock_lower_row_out => s_locks_lower_out(8,40),
			lock_lower_row_in  => s_locks_lower_in(8,40),
			in1                => s_in1(8,40),
			in2                => s_in2(8,40),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(40)
		);
	s_in1(8,40)            <= s_out1(9,40);
	s_in2(8,40)            <= s_out2(9,41);
	s_locks_lower_in(8,40) <= s_locks_lower_out(9,40);

		normal_cell_8_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,41),
			fetch              => s_fetch(8,41),
			data_in            => s_data_in(8,41),
			data_out           => s_data_out(8,41),
			out1               => s_out1(8,41),
			out2               => s_out2(8,41),
			lock_lower_row_out => s_locks_lower_out(8,41),
			lock_lower_row_in  => s_locks_lower_in(8,41),
			in1                => s_in1(8,41),
			in2                => s_in2(8,41),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(41)
		);
	s_in1(8,41)            <= s_out1(9,41);
	s_in2(8,41)            <= s_out2(9,42);
	s_locks_lower_in(8,41) <= s_locks_lower_out(9,41);

		normal_cell_8_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,42),
			fetch              => s_fetch(8,42),
			data_in            => s_data_in(8,42),
			data_out           => s_data_out(8,42),
			out1               => s_out1(8,42),
			out2               => s_out2(8,42),
			lock_lower_row_out => s_locks_lower_out(8,42),
			lock_lower_row_in  => s_locks_lower_in(8,42),
			in1                => s_in1(8,42),
			in2                => s_in2(8,42),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(42)
		);
	s_in1(8,42)            <= s_out1(9,42);
	s_in2(8,42)            <= s_out2(9,43);
	s_locks_lower_in(8,42) <= s_locks_lower_out(9,42);

		normal_cell_8_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,43),
			fetch              => s_fetch(8,43),
			data_in            => s_data_in(8,43),
			data_out           => s_data_out(8,43),
			out1               => s_out1(8,43),
			out2               => s_out2(8,43),
			lock_lower_row_out => s_locks_lower_out(8,43),
			lock_lower_row_in  => s_locks_lower_in(8,43),
			in1                => s_in1(8,43),
			in2                => s_in2(8,43),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(43)
		);
	s_in1(8,43)            <= s_out1(9,43);
	s_in2(8,43)            <= s_out2(9,44);
	s_locks_lower_in(8,43) <= s_locks_lower_out(9,43);

		normal_cell_8_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,44),
			fetch              => s_fetch(8,44),
			data_in            => s_data_in(8,44),
			data_out           => s_data_out(8,44),
			out1               => s_out1(8,44),
			out2               => s_out2(8,44),
			lock_lower_row_out => s_locks_lower_out(8,44),
			lock_lower_row_in  => s_locks_lower_in(8,44),
			in1                => s_in1(8,44),
			in2                => s_in2(8,44),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(44)
		);
	s_in1(8,44)            <= s_out1(9,44);
	s_in2(8,44)            <= s_out2(9,45);
	s_locks_lower_in(8,44) <= s_locks_lower_out(9,44);

		normal_cell_8_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,45),
			fetch              => s_fetch(8,45),
			data_in            => s_data_in(8,45),
			data_out           => s_data_out(8,45),
			out1               => s_out1(8,45),
			out2               => s_out2(8,45),
			lock_lower_row_out => s_locks_lower_out(8,45),
			lock_lower_row_in  => s_locks_lower_in(8,45),
			in1                => s_in1(8,45),
			in2                => s_in2(8,45),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(45)
		);
	s_in1(8,45)            <= s_out1(9,45);
	s_in2(8,45)            <= s_out2(9,46);
	s_locks_lower_in(8,45) <= s_locks_lower_out(9,45);

		normal_cell_8_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,46),
			fetch              => s_fetch(8,46),
			data_in            => s_data_in(8,46),
			data_out           => s_data_out(8,46),
			out1               => s_out1(8,46),
			out2               => s_out2(8,46),
			lock_lower_row_out => s_locks_lower_out(8,46),
			lock_lower_row_in  => s_locks_lower_in(8,46),
			in1                => s_in1(8,46),
			in2                => s_in2(8,46),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(46)
		);
	s_in1(8,46)            <= s_out1(9,46);
	s_in2(8,46)            <= s_out2(9,47);
	s_locks_lower_in(8,46) <= s_locks_lower_out(9,46);

		normal_cell_8_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,47),
			fetch              => s_fetch(8,47),
			data_in            => s_data_in(8,47),
			data_out           => s_data_out(8,47),
			out1               => s_out1(8,47),
			out2               => s_out2(8,47),
			lock_lower_row_out => s_locks_lower_out(8,47),
			lock_lower_row_in  => s_locks_lower_in(8,47),
			in1                => s_in1(8,47),
			in2                => s_in2(8,47),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(47)
		);
	s_in1(8,47)            <= s_out1(9,47);
	s_in2(8,47)            <= s_out2(9,48);
	s_locks_lower_in(8,47) <= s_locks_lower_out(9,47);

		normal_cell_8_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,48),
			fetch              => s_fetch(8,48),
			data_in            => s_data_in(8,48),
			data_out           => s_data_out(8,48),
			out1               => s_out1(8,48),
			out2               => s_out2(8,48),
			lock_lower_row_out => s_locks_lower_out(8,48),
			lock_lower_row_in  => s_locks_lower_in(8,48),
			in1                => s_in1(8,48),
			in2                => s_in2(8,48),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(48)
		);
	s_in1(8,48)            <= s_out1(9,48);
	s_in2(8,48)            <= s_out2(9,49);
	s_locks_lower_in(8,48) <= s_locks_lower_out(9,48);

		normal_cell_8_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,49),
			fetch              => s_fetch(8,49),
			data_in            => s_data_in(8,49),
			data_out           => s_data_out(8,49),
			out1               => s_out1(8,49),
			out2               => s_out2(8,49),
			lock_lower_row_out => s_locks_lower_out(8,49),
			lock_lower_row_in  => s_locks_lower_in(8,49),
			in1                => s_in1(8,49),
			in2                => s_in2(8,49),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(49)
		);
	s_in1(8,49)            <= s_out1(9,49);
	s_in2(8,49)            <= s_out2(9,50);
	s_locks_lower_in(8,49) <= s_locks_lower_out(9,49);

		normal_cell_8_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,50),
			fetch              => s_fetch(8,50),
			data_in            => s_data_in(8,50),
			data_out           => s_data_out(8,50),
			out1               => s_out1(8,50),
			out2               => s_out2(8,50),
			lock_lower_row_out => s_locks_lower_out(8,50),
			lock_lower_row_in  => s_locks_lower_in(8,50),
			in1                => s_in1(8,50),
			in2                => s_in2(8,50),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(50)
		);
	s_in1(8,50)            <= s_out1(9,50);
	s_in2(8,50)            <= s_out2(9,51);
	s_locks_lower_in(8,50) <= s_locks_lower_out(9,50);

		normal_cell_8_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,51),
			fetch              => s_fetch(8,51),
			data_in            => s_data_in(8,51),
			data_out           => s_data_out(8,51),
			out1               => s_out1(8,51),
			out2               => s_out2(8,51),
			lock_lower_row_out => s_locks_lower_out(8,51),
			lock_lower_row_in  => s_locks_lower_in(8,51),
			in1                => s_in1(8,51),
			in2                => s_in2(8,51),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(51)
		);
	s_in1(8,51)            <= s_out1(9,51);
	s_in2(8,51)            <= s_out2(9,52);
	s_locks_lower_in(8,51) <= s_locks_lower_out(9,51);

		normal_cell_8_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,52),
			fetch              => s_fetch(8,52),
			data_in            => s_data_in(8,52),
			data_out           => s_data_out(8,52),
			out1               => s_out1(8,52),
			out2               => s_out2(8,52),
			lock_lower_row_out => s_locks_lower_out(8,52),
			lock_lower_row_in  => s_locks_lower_in(8,52),
			in1                => s_in1(8,52),
			in2                => s_in2(8,52),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(52)
		);
	s_in1(8,52)            <= s_out1(9,52);
	s_in2(8,52)            <= s_out2(9,53);
	s_locks_lower_in(8,52) <= s_locks_lower_out(9,52);

		normal_cell_8_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,53),
			fetch              => s_fetch(8,53),
			data_in            => s_data_in(8,53),
			data_out           => s_data_out(8,53),
			out1               => s_out1(8,53),
			out2               => s_out2(8,53),
			lock_lower_row_out => s_locks_lower_out(8,53),
			lock_lower_row_in  => s_locks_lower_in(8,53),
			in1                => s_in1(8,53),
			in2                => s_in2(8,53),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(53)
		);
	s_in1(8,53)            <= s_out1(9,53);
	s_in2(8,53)            <= s_out2(9,54);
	s_locks_lower_in(8,53) <= s_locks_lower_out(9,53);

		normal_cell_8_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,54),
			fetch              => s_fetch(8,54),
			data_in            => s_data_in(8,54),
			data_out           => s_data_out(8,54),
			out1               => s_out1(8,54),
			out2               => s_out2(8,54),
			lock_lower_row_out => s_locks_lower_out(8,54),
			lock_lower_row_in  => s_locks_lower_in(8,54),
			in1                => s_in1(8,54),
			in2                => s_in2(8,54),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(54)
		);
	s_in1(8,54)            <= s_out1(9,54);
	s_in2(8,54)            <= s_out2(9,55);
	s_locks_lower_in(8,54) <= s_locks_lower_out(9,54);

		normal_cell_8_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,55),
			fetch              => s_fetch(8,55),
			data_in            => s_data_in(8,55),
			data_out           => s_data_out(8,55),
			out1               => s_out1(8,55),
			out2               => s_out2(8,55),
			lock_lower_row_out => s_locks_lower_out(8,55),
			lock_lower_row_in  => s_locks_lower_in(8,55),
			in1                => s_in1(8,55),
			in2                => s_in2(8,55),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(55)
		);
	s_in1(8,55)            <= s_out1(9,55);
	s_in2(8,55)            <= s_out2(9,56);
	s_locks_lower_in(8,55) <= s_locks_lower_out(9,55);

		normal_cell_8_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,56),
			fetch              => s_fetch(8,56),
			data_in            => s_data_in(8,56),
			data_out           => s_data_out(8,56),
			out1               => s_out1(8,56),
			out2               => s_out2(8,56),
			lock_lower_row_out => s_locks_lower_out(8,56),
			lock_lower_row_in  => s_locks_lower_in(8,56),
			in1                => s_in1(8,56),
			in2                => s_in2(8,56),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(56)
		);
	s_in1(8,56)            <= s_out1(9,56);
	s_in2(8,56)            <= s_out2(9,57);
	s_locks_lower_in(8,56) <= s_locks_lower_out(9,56);

		normal_cell_8_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,57),
			fetch              => s_fetch(8,57),
			data_in            => s_data_in(8,57),
			data_out           => s_data_out(8,57),
			out1               => s_out1(8,57),
			out2               => s_out2(8,57),
			lock_lower_row_out => s_locks_lower_out(8,57),
			lock_lower_row_in  => s_locks_lower_in(8,57),
			in1                => s_in1(8,57),
			in2                => s_in2(8,57),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(57)
		);
	s_in1(8,57)            <= s_out1(9,57);
	s_in2(8,57)            <= s_out2(9,58);
	s_locks_lower_in(8,57) <= s_locks_lower_out(9,57);

		normal_cell_8_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,58),
			fetch              => s_fetch(8,58),
			data_in            => s_data_in(8,58),
			data_out           => s_data_out(8,58),
			out1               => s_out1(8,58),
			out2               => s_out2(8,58),
			lock_lower_row_out => s_locks_lower_out(8,58),
			lock_lower_row_in  => s_locks_lower_in(8,58),
			in1                => s_in1(8,58),
			in2                => s_in2(8,58),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(58)
		);
	s_in1(8,58)            <= s_out1(9,58);
	s_in2(8,58)            <= s_out2(9,59);
	s_locks_lower_in(8,58) <= s_locks_lower_out(9,58);

		normal_cell_8_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,59),
			fetch              => s_fetch(8,59),
			data_in            => s_data_in(8,59),
			data_out           => s_data_out(8,59),
			out1               => s_out1(8,59),
			out2               => s_out2(8,59),
			lock_lower_row_out => s_locks_lower_out(8,59),
			lock_lower_row_in  => s_locks_lower_in(8,59),
			in1                => s_in1(8,59),
			in2                => s_in2(8,59),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(59)
		);
	s_in1(8,59)            <= s_out1(9,59);
	s_in2(8,59)            <= s_out2(9,60);
	s_locks_lower_in(8,59) <= s_locks_lower_out(9,59);

		last_col_cell_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(8,60),
			fetch              => s_fetch(8,60),
			data_in            => s_data_in(8,60),
			data_out           => s_data_out(8,60),
			out1               => s_out1(8,60),
			out2               => s_out2(8,60),
			lock_lower_row_out => s_locks_lower_out(8,60),
			lock_lower_row_in  => s_locks_lower_in(8,60),
			in1                => s_in1(8,60),
			in2                => (others => '0'),
			lock_row           => s_locks(8),
			piv_found          => s_piv_found,
			row_data           => s_row_data(8),
			col_data           => s_col_data(60)
		);
	s_in1(8,60)            <= s_out1(9,60);
	s_locks_lower_in(8,60) <= s_locks_lower_out(9,60);

		normal_cell_9_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,1),
			fetch              => s_fetch(9,1),
			data_in            => s_data_in(9,1),
			data_out           => s_data_out(9,1),
			out1               => s_out1(9,1),
			out2               => s_out2(9,1),
			lock_lower_row_out => s_locks_lower_out(9,1),
			lock_lower_row_in  => s_locks_lower_in(9,1),
			in1                => s_in1(9,1),
			in2                => s_in2(9,1),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(1)
		);
	s_in1(9,1)            <= s_out1(10,1);
	s_in2(9,1)            <= s_out2(10,2);
	s_locks_lower_in(9,1) <= s_locks_lower_out(10,1);

		normal_cell_9_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,2),
			fetch              => s_fetch(9,2),
			data_in            => s_data_in(9,2),
			data_out           => s_data_out(9,2),
			out1               => s_out1(9,2),
			out2               => s_out2(9,2),
			lock_lower_row_out => s_locks_lower_out(9,2),
			lock_lower_row_in  => s_locks_lower_in(9,2),
			in1                => s_in1(9,2),
			in2                => s_in2(9,2),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(2)
		);
	s_in1(9,2)            <= s_out1(10,2);
	s_in2(9,2)            <= s_out2(10,3);
	s_locks_lower_in(9,2) <= s_locks_lower_out(10,2);

		normal_cell_9_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,3),
			fetch              => s_fetch(9,3),
			data_in            => s_data_in(9,3),
			data_out           => s_data_out(9,3),
			out1               => s_out1(9,3),
			out2               => s_out2(9,3),
			lock_lower_row_out => s_locks_lower_out(9,3),
			lock_lower_row_in  => s_locks_lower_in(9,3),
			in1                => s_in1(9,3),
			in2                => s_in2(9,3),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(3)
		);
	s_in1(9,3)            <= s_out1(10,3);
	s_in2(9,3)            <= s_out2(10,4);
	s_locks_lower_in(9,3) <= s_locks_lower_out(10,3);

		normal_cell_9_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,4),
			fetch              => s_fetch(9,4),
			data_in            => s_data_in(9,4),
			data_out           => s_data_out(9,4),
			out1               => s_out1(9,4),
			out2               => s_out2(9,4),
			lock_lower_row_out => s_locks_lower_out(9,4),
			lock_lower_row_in  => s_locks_lower_in(9,4),
			in1                => s_in1(9,4),
			in2                => s_in2(9,4),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(4)
		);
	s_in1(9,4)            <= s_out1(10,4);
	s_in2(9,4)            <= s_out2(10,5);
	s_locks_lower_in(9,4) <= s_locks_lower_out(10,4);

		normal_cell_9_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,5),
			fetch              => s_fetch(9,5),
			data_in            => s_data_in(9,5),
			data_out           => s_data_out(9,5),
			out1               => s_out1(9,5),
			out2               => s_out2(9,5),
			lock_lower_row_out => s_locks_lower_out(9,5),
			lock_lower_row_in  => s_locks_lower_in(9,5),
			in1                => s_in1(9,5),
			in2                => s_in2(9,5),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(5)
		);
	s_in1(9,5)            <= s_out1(10,5);
	s_in2(9,5)            <= s_out2(10,6);
	s_locks_lower_in(9,5) <= s_locks_lower_out(10,5);

		normal_cell_9_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,6),
			fetch              => s_fetch(9,6),
			data_in            => s_data_in(9,6),
			data_out           => s_data_out(9,6),
			out1               => s_out1(9,6),
			out2               => s_out2(9,6),
			lock_lower_row_out => s_locks_lower_out(9,6),
			lock_lower_row_in  => s_locks_lower_in(9,6),
			in1                => s_in1(9,6),
			in2                => s_in2(9,6),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(6)
		);
	s_in1(9,6)            <= s_out1(10,6);
	s_in2(9,6)            <= s_out2(10,7);
	s_locks_lower_in(9,6) <= s_locks_lower_out(10,6);

		normal_cell_9_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,7),
			fetch              => s_fetch(9,7),
			data_in            => s_data_in(9,7),
			data_out           => s_data_out(9,7),
			out1               => s_out1(9,7),
			out2               => s_out2(9,7),
			lock_lower_row_out => s_locks_lower_out(9,7),
			lock_lower_row_in  => s_locks_lower_in(9,7),
			in1                => s_in1(9,7),
			in2                => s_in2(9,7),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(7)
		);
	s_in1(9,7)            <= s_out1(10,7);
	s_in2(9,7)            <= s_out2(10,8);
	s_locks_lower_in(9,7) <= s_locks_lower_out(10,7);

		normal_cell_9_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,8),
			fetch              => s_fetch(9,8),
			data_in            => s_data_in(9,8),
			data_out           => s_data_out(9,8),
			out1               => s_out1(9,8),
			out2               => s_out2(9,8),
			lock_lower_row_out => s_locks_lower_out(9,8),
			lock_lower_row_in  => s_locks_lower_in(9,8),
			in1                => s_in1(9,8),
			in2                => s_in2(9,8),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(8)
		);
	s_in1(9,8)            <= s_out1(10,8);
	s_in2(9,8)            <= s_out2(10,9);
	s_locks_lower_in(9,8) <= s_locks_lower_out(10,8);

		normal_cell_9_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,9),
			fetch              => s_fetch(9,9),
			data_in            => s_data_in(9,9),
			data_out           => s_data_out(9,9),
			out1               => s_out1(9,9),
			out2               => s_out2(9,9),
			lock_lower_row_out => s_locks_lower_out(9,9),
			lock_lower_row_in  => s_locks_lower_in(9,9),
			in1                => s_in1(9,9),
			in2                => s_in2(9,9),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(9)
		);
	s_in1(9,9)            <= s_out1(10,9);
	s_in2(9,9)            <= s_out2(10,10);
	s_locks_lower_in(9,9) <= s_locks_lower_out(10,9);

		normal_cell_9_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,10),
			fetch              => s_fetch(9,10),
			data_in            => s_data_in(9,10),
			data_out           => s_data_out(9,10),
			out1               => s_out1(9,10),
			out2               => s_out2(9,10),
			lock_lower_row_out => s_locks_lower_out(9,10),
			lock_lower_row_in  => s_locks_lower_in(9,10),
			in1                => s_in1(9,10),
			in2                => s_in2(9,10),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(10)
		);
	s_in1(9,10)            <= s_out1(10,10);
	s_in2(9,10)            <= s_out2(10,11);
	s_locks_lower_in(9,10) <= s_locks_lower_out(10,10);

		normal_cell_9_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,11),
			fetch              => s_fetch(9,11),
			data_in            => s_data_in(9,11),
			data_out           => s_data_out(9,11),
			out1               => s_out1(9,11),
			out2               => s_out2(9,11),
			lock_lower_row_out => s_locks_lower_out(9,11),
			lock_lower_row_in  => s_locks_lower_in(9,11),
			in1                => s_in1(9,11),
			in2                => s_in2(9,11),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(11)
		);
	s_in1(9,11)            <= s_out1(10,11);
	s_in2(9,11)            <= s_out2(10,12);
	s_locks_lower_in(9,11) <= s_locks_lower_out(10,11);

		normal_cell_9_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,12),
			fetch              => s_fetch(9,12),
			data_in            => s_data_in(9,12),
			data_out           => s_data_out(9,12),
			out1               => s_out1(9,12),
			out2               => s_out2(9,12),
			lock_lower_row_out => s_locks_lower_out(9,12),
			lock_lower_row_in  => s_locks_lower_in(9,12),
			in1                => s_in1(9,12),
			in2                => s_in2(9,12),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(12)
		);
	s_in1(9,12)            <= s_out1(10,12);
	s_in2(9,12)            <= s_out2(10,13);
	s_locks_lower_in(9,12) <= s_locks_lower_out(10,12);

		normal_cell_9_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,13),
			fetch              => s_fetch(9,13),
			data_in            => s_data_in(9,13),
			data_out           => s_data_out(9,13),
			out1               => s_out1(9,13),
			out2               => s_out2(9,13),
			lock_lower_row_out => s_locks_lower_out(9,13),
			lock_lower_row_in  => s_locks_lower_in(9,13),
			in1                => s_in1(9,13),
			in2                => s_in2(9,13),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(13)
		);
	s_in1(9,13)            <= s_out1(10,13);
	s_in2(9,13)            <= s_out2(10,14);
	s_locks_lower_in(9,13) <= s_locks_lower_out(10,13);

		normal_cell_9_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,14),
			fetch              => s_fetch(9,14),
			data_in            => s_data_in(9,14),
			data_out           => s_data_out(9,14),
			out1               => s_out1(9,14),
			out2               => s_out2(9,14),
			lock_lower_row_out => s_locks_lower_out(9,14),
			lock_lower_row_in  => s_locks_lower_in(9,14),
			in1                => s_in1(9,14),
			in2                => s_in2(9,14),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(14)
		);
	s_in1(9,14)            <= s_out1(10,14);
	s_in2(9,14)            <= s_out2(10,15);
	s_locks_lower_in(9,14) <= s_locks_lower_out(10,14);

		normal_cell_9_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,15),
			fetch              => s_fetch(9,15),
			data_in            => s_data_in(9,15),
			data_out           => s_data_out(9,15),
			out1               => s_out1(9,15),
			out2               => s_out2(9,15),
			lock_lower_row_out => s_locks_lower_out(9,15),
			lock_lower_row_in  => s_locks_lower_in(9,15),
			in1                => s_in1(9,15),
			in2                => s_in2(9,15),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(15)
		);
	s_in1(9,15)            <= s_out1(10,15);
	s_in2(9,15)            <= s_out2(10,16);
	s_locks_lower_in(9,15) <= s_locks_lower_out(10,15);

		normal_cell_9_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,16),
			fetch              => s_fetch(9,16),
			data_in            => s_data_in(9,16),
			data_out           => s_data_out(9,16),
			out1               => s_out1(9,16),
			out2               => s_out2(9,16),
			lock_lower_row_out => s_locks_lower_out(9,16),
			lock_lower_row_in  => s_locks_lower_in(9,16),
			in1                => s_in1(9,16),
			in2                => s_in2(9,16),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(16)
		);
	s_in1(9,16)            <= s_out1(10,16);
	s_in2(9,16)            <= s_out2(10,17);
	s_locks_lower_in(9,16) <= s_locks_lower_out(10,16);

		normal_cell_9_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,17),
			fetch              => s_fetch(9,17),
			data_in            => s_data_in(9,17),
			data_out           => s_data_out(9,17),
			out1               => s_out1(9,17),
			out2               => s_out2(9,17),
			lock_lower_row_out => s_locks_lower_out(9,17),
			lock_lower_row_in  => s_locks_lower_in(9,17),
			in1                => s_in1(9,17),
			in2                => s_in2(9,17),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(17)
		);
	s_in1(9,17)            <= s_out1(10,17);
	s_in2(9,17)            <= s_out2(10,18);
	s_locks_lower_in(9,17) <= s_locks_lower_out(10,17);

		normal_cell_9_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,18),
			fetch              => s_fetch(9,18),
			data_in            => s_data_in(9,18),
			data_out           => s_data_out(9,18),
			out1               => s_out1(9,18),
			out2               => s_out2(9,18),
			lock_lower_row_out => s_locks_lower_out(9,18),
			lock_lower_row_in  => s_locks_lower_in(9,18),
			in1                => s_in1(9,18),
			in2                => s_in2(9,18),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(18)
		);
	s_in1(9,18)            <= s_out1(10,18);
	s_in2(9,18)            <= s_out2(10,19);
	s_locks_lower_in(9,18) <= s_locks_lower_out(10,18);

		normal_cell_9_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,19),
			fetch              => s_fetch(9,19),
			data_in            => s_data_in(9,19),
			data_out           => s_data_out(9,19),
			out1               => s_out1(9,19),
			out2               => s_out2(9,19),
			lock_lower_row_out => s_locks_lower_out(9,19),
			lock_lower_row_in  => s_locks_lower_in(9,19),
			in1                => s_in1(9,19),
			in2                => s_in2(9,19),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(19)
		);
	s_in1(9,19)            <= s_out1(10,19);
	s_in2(9,19)            <= s_out2(10,20);
	s_locks_lower_in(9,19) <= s_locks_lower_out(10,19);

		normal_cell_9_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,20),
			fetch              => s_fetch(9,20),
			data_in            => s_data_in(9,20),
			data_out           => s_data_out(9,20),
			out1               => s_out1(9,20),
			out2               => s_out2(9,20),
			lock_lower_row_out => s_locks_lower_out(9,20),
			lock_lower_row_in  => s_locks_lower_in(9,20),
			in1                => s_in1(9,20),
			in2                => s_in2(9,20),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(20)
		);
	s_in1(9,20)            <= s_out1(10,20);
	s_in2(9,20)            <= s_out2(10,21);
	s_locks_lower_in(9,20) <= s_locks_lower_out(10,20);

		normal_cell_9_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,21),
			fetch              => s_fetch(9,21),
			data_in            => s_data_in(9,21),
			data_out           => s_data_out(9,21),
			out1               => s_out1(9,21),
			out2               => s_out2(9,21),
			lock_lower_row_out => s_locks_lower_out(9,21),
			lock_lower_row_in  => s_locks_lower_in(9,21),
			in1                => s_in1(9,21),
			in2                => s_in2(9,21),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(21)
		);
	s_in1(9,21)            <= s_out1(10,21);
	s_in2(9,21)            <= s_out2(10,22);
	s_locks_lower_in(9,21) <= s_locks_lower_out(10,21);

		normal_cell_9_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,22),
			fetch              => s_fetch(9,22),
			data_in            => s_data_in(9,22),
			data_out           => s_data_out(9,22),
			out1               => s_out1(9,22),
			out2               => s_out2(9,22),
			lock_lower_row_out => s_locks_lower_out(9,22),
			lock_lower_row_in  => s_locks_lower_in(9,22),
			in1                => s_in1(9,22),
			in2                => s_in2(9,22),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(22)
		);
	s_in1(9,22)            <= s_out1(10,22);
	s_in2(9,22)            <= s_out2(10,23);
	s_locks_lower_in(9,22) <= s_locks_lower_out(10,22);

		normal_cell_9_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,23),
			fetch              => s_fetch(9,23),
			data_in            => s_data_in(9,23),
			data_out           => s_data_out(9,23),
			out1               => s_out1(9,23),
			out2               => s_out2(9,23),
			lock_lower_row_out => s_locks_lower_out(9,23),
			lock_lower_row_in  => s_locks_lower_in(9,23),
			in1                => s_in1(9,23),
			in2                => s_in2(9,23),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(23)
		);
	s_in1(9,23)            <= s_out1(10,23);
	s_in2(9,23)            <= s_out2(10,24);
	s_locks_lower_in(9,23) <= s_locks_lower_out(10,23);

		normal_cell_9_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,24),
			fetch              => s_fetch(9,24),
			data_in            => s_data_in(9,24),
			data_out           => s_data_out(9,24),
			out1               => s_out1(9,24),
			out2               => s_out2(9,24),
			lock_lower_row_out => s_locks_lower_out(9,24),
			lock_lower_row_in  => s_locks_lower_in(9,24),
			in1                => s_in1(9,24),
			in2                => s_in2(9,24),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(24)
		);
	s_in1(9,24)            <= s_out1(10,24);
	s_in2(9,24)            <= s_out2(10,25);
	s_locks_lower_in(9,24) <= s_locks_lower_out(10,24);

		normal_cell_9_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,25),
			fetch              => s_fetch(9,25),
			data_in            => s_data_in(9,25),
			data_out           => s_data_out(9,25),
			out1               => s_out1(9,25),
			out2               => s_out2(9,25),
			lock_lower_row_out => s_locks_lower_out(9,25),
			lock_lower_row_in  => s_locks_lower_in(9,25),
			in1                => s_in1(9,25),
			in2                => s_in2(9,25),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(25)
		);
	s_in1(9,25)            <= s_out1(10,25);
	s_in2(9,25)            <= s_out2(10,26);
	s_locks_lower_in(9,25) <= s_locks_lower_out(10,25);

		normal_cell_9_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,26),
			fetch              => s_fetch(9,26),
			data_in            => s_data_in(9,26),
			data_out           => s_data_out(9,26),
			out1               => s_out1(9,26),
			out2               => s_out2(9,26),
			lock_lower_row_out => s_locks_lower_out(9,26),
			lock_lower_row_in  => s_locks_lower_in(9,26),
			in1                => s_in1(9,26),
			in2                => s_in2(9,26),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(26)
		);
	s_in1(9,26)            <= s_out1(10,26);
	s_in2(9,26)            <= s_out2(10,27);
	s_locks_lower_in(9,26) <= s_locks_lower_out(10,26);

		normal_cell_9_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,27),
			fetch              => s_fetch(9,27),
			data_in            => s_data_in(9,27),
			data_out           => s_data_out(9,27),
			out1               => s_out1(9,27),
			out2               => s_out2(9,27),
			lock_lower_row_out => s_locks_lower_out(9,27),
			lock_lower_row_in  => s_locks_lower_in(9,27),
			in1                => s_in1(9,27),
			in2                => s_in2(9,27),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(27)
		);
	s_in1(9,27)            <= s_out1(10,27);
	s_in2(9,27)            <= s_out2(10,28);
	s_locks_lower_in(9,27) <= s_locks_lower_out(10,27);

		normal_cell_9_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,28),
			fetch              => s_fetch(9,28),
			data_in            => s_data_in(9,28),
			data_out           => s_data_out(9,28),
			out1               => s_out1(9,28),
			out2               => s_out2(9,28),
			lock_lower_row_out => s_locks_lower_out(9,28),
			lock_lower_row_in  => s_locks_lower_in(9,28),
			in1                => s_in1(9,28),
			in2                => s_in2(9,28),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(28)
		);
	s_in1(9,28)            <= s_out1(10,28);
	s_in2(9,28)            <= s_out2(10,29);
	s_locks_lower_in(9,28) <= s_locks_lower_out(10,28);

		normal_cell_9_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,29),
			fetch              => s_fetch(9,29),
			data_in            => s_data_in(9,29),
			data_out           => s_data_out(9,29),
			out1               => s_out1(9,29),
			out2               => s_out2(9,29),
			lock_lower_row_out => s_locks_lower_out(9,29),
			lock_lower_row_in  => s_locks_lower_in(9,29),
			in1                => s_in1(9,29),
			in2                => s_in2(9,29),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(29)
		);
	s_in1(9,29)            <= s_out1(10,29);
	s_in2(9,29)            <= s_out2(10,30);
	s_locks_lower_in(9,29) <= s_locks_lower_out(10,29);

		normal_cell_9_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,30),
			fetch              => s_fetch(9,30),
			data_in            => s_data_in(9,30),
			data_out           => s_data_out(9,30),
			out1               => s_out1(9,30),
			out2               => s_out2(9,30),
			lock_lower_row_out => s_locks_lower_out(9,30),
			lock_lower_row_in  => s_locks_lower_in(9,30),
			in1                => s_in1(9,30),
			in2                => s_in2(9,30),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(30)
		);
	s_in1(9,30)            <= s_out1(10,30);
	s_in2(9,30)            <= s_out2(10,31);
	s_locks_lower_in(9,30) <= s_locks_lower_out(10,30);

		normal_cell_9_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,31),
			fetch              => s_fetch(9,31),
			data_in            => s_data_in(9,31),
			data_out           => s_data_out(9,31),
			out1               => s_out1(9,31),
			out2               => s_out2(9,31),
			lock_lower_row_out => s_locks_lower_out(9,31),
			lock_lower_row_in  => s_locks_lower_in(9,31),
			in1                => s_in1(9,31),
			in2                => s_in2(9,31),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(31)
		);
	s_in1(9,31)            <= s_out1(10,31);
	s_in2(9,31)            <= s_out2(10,32);
	s_locks_lower_in(9,31) <= s_locks_lower_out(10,31);

		normal_cell_9_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,32),
			fetch              => s_fetch(9,32),
			data_in            => s_data_in(9,32),
			data_out           => s_data_out(9,32),
			out1               => s_out1(9,32),
			out2               => s_out2(9,32),
			lock_lower_row_out => s_locks_lower_out(9,32),
			lock_lower_row_in  => s_locks_lower_in(9,32),
			in1                => s_in1(9,32),
			in2                => s_in2(9,32),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(32)
		);
	s_in1(9,32)            <= s_out1(10,32);
	s_in2(9,32)            <= s_out2(10,33);
	s_locks_lower_in(9,32) <= s_locks_lower_out(10,32);

		normal_cell_9_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,33),
			fetch              => s_fetch(9,33),
			data_in            => s_data_in(9,33),
			data_out           => s_data_out(9,33),
			out1               => s_out1(9,33),
			out2               => s_out2(9,33),
			lock_lower_row_out => s_locks_lower_out(9,33),
			lock_lower_row_in  => s_locks_lower_in(9,33),
			in1                => s_in1(9,33),
			in2                => s_in2(9,33),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(33)
		);
	s_in1(9,33)            <= s_out1(10,33);
	s_in2(9,33)            <= s_out2(10,34);
	s_locks_lower_in(9,33) <= s_locks_lower_out(10,33);

		normal_cell_9_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,34),
			fetch              => s_fetch(9,34),
			data_in            => s_data_in(9,34),
			data_out           => s_data_out(9,34),
			out1               => s_out1(9,34),
			out2               => s_out2(9,34),
			lock_lower_row_out => s_locks_lower_out(9,34),
			lock_lower_row_in  => s_locks_lower_in(9,34),
			in1                => s_in1(9,34),
			in2                => s_in2(9,34),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(34)
		);
	s_in1(9,34)            <= s_out1(10,34);
	s_in2(9,34)            <= s_out2(10,35);
	s_locks_lower_in(9,34) <= s_locks_lower_out(10,34);

		normal_cell_9_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,35),
			fetch              => s_fetch(9,35),
			data_in            => s_data_in(9,35),
			data_out           => s_data_out(9,35),
			out1               => s_out1(9,35),
			out2               => s_out2(9,35),
			lock_lower_row_out => s_locks_lower_out(9,35),
			lock_lower_row_in  => s_locks_lower_in(9,35),
			in1                => s_in1(9,35),
			in2                => s_in2(9,35),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(35)
		);
	s_in1(9,35)            <= s_out1(10,35);
	s_in2(9,35)            <= s_out2(10,36);
	s_locks_lower_in(9,35) <= s_locks_lower_out(10,35);

		normal_cell_9_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,36),
			fetch              => s_fetch(9,36),
			data_in            => s_data_in(9,36),
			data_out           => s_data_out(9,36),
			out1               => s_out1(9,36),
			out2               => s_out2(9,36),
			lock_lower_row_out => s_locks_lower_out(9,36),
			lock_lower_row_in  => s_locks_lower_in(9,36),
			in1                => s_in1(9,36),
			in2                => s_in2(9,36),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(36)
		);
	s_in1(9,36)            <= s_out1(10,36);
	s_in2(9,36)            <= s_out2(10,37);
	s_locks_lower_in(9,36) <= s_locks_lower_out(10,36);

		normal_cell_9_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,37),
			fetch              => s_fetch(9,37),
			data_in            => s_data_in(9,37),
			data_out           => s_data_out(9,37),
			out1               => s_out1(9,37),
			out2               => s_out2(9,37),
			lock_lower_row_out => s_locks_lower_out(9,37),
			lock_lower_row_in  => s_locks_lower_in(9,37),
			in1                => s_in1(9,37),
			in2                => s_in2(9,37),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(37)
		);
	s_in1(9,37)            <= s_out1(10,37);
	s_in2(9,37)            <= s_out2(10,38);
	s_locks_lower_in(9,37) <= s_locks_lower_out(10,37);

		normal_cell_9_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,38),
			fetch              => s_fetch(9,38),
			data_in            => s_data_in(9,38),
			data_out           => s_data_out(9,38),
			out1               => s_out1(9,38),
			out2               => s_out2(9,38),
			lock_lower_row_out => s_locks_lower_out(9,38),
			lock_lower_row_in  => s_locks_lower_in(9,38),
			in1                => s_in1(9,38),
			in2                => s_in2(9,38),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(38)
		);
	s_in1(9,38)            <= s_out1(10,38);
	s_in2(9,38)            <= s_out2(10,39);
	s_locks_lower_in(9,38) <= s_locks_lower_out(10,38);

		normal_cell_9_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,39),
			fetch              => s_fetch(9,39),
			data_in            => s_data_in(9,39),
			data_out           => s_data_out(9,39),
			out1               => s_out1(9,39),
			out2               => s_out2(9,39),
			lock_lower_row_out => s_locks_lower_out(9,39),
			lock_lower_row_in  => s_locks_lower_in(9,39),
			in1                => s_in1(9,39),
			in2                => s_in2(9,39),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(39)
		);
	s_in1(9,39)            <= s_out1(10,39);
	s_in2(9,39)            <= s_out2(10,40);
	s_locks_lower_in(9,39) <= s_locks_lower_out(10,39);

		normal_cell_9_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,40),
			fetch              => s_fetch(9,40),
			data_in            => s_data_in(9,40),
			data_out           => s_data_out(9,40),
			out1               => s_out1(9,40),
			out2               => s_out2(9,40),
			lock_lower_row_out => s_locks_lower_out(9,40),
			lock_lower_row_in  => s_locks_lower_in(9,40),
			in1                => s_in1(9,40),
			in2                => s_in2(9,40),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(40)
		);
	s_in1(9,40)            <= s_out1(10,40);
	s_in2(9,40)            <= s_out2(10,41);
	s_locks_lower_in(9,40) <= s_locks_lower_out(10,40);

		normal_cell_9_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,41),
			fetch              => s_fetch(9,41),
			data_in            => s_data_in(9,41),
			data_out           => s_data_out(9,41),
			out1               => s_out1(9,41),
			out2               => s_out2(9,41),
			lock_lower_row_out => s_locks_lower_out(9,41),
			lock_lower_row_in  => s_locks_lower_in(9,41),
			in1                => s_in1(9,41),
			in2                => s_in2(9,41),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(41)
		);
	s_in1(9,41)            <= s_out1(10,41);
	s_in2(9,41)            <= s_out2(10,42);
	s_locks_lower_in(9,41) <= s_locks_lower_out(10,41);

		normal_cell_9_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,42),
			fetch              => s_fetch(9,42),
			data_in            => s_data_in(9,42),
			data_out           => s_data_out(9,42),
			out1               => s_out1(9,42),
			out2               => s_out2(9,42),
			lock_lower_row_out => s_locks_lower_out(9,42),
			lock_lower_row_in  => s_locks_lower_in(9,42),
			in1                => s_in1(9,42),
			in2                => s_in2(9,42),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(42)
		);
	s_in1(9,42)            <= s_out1(10,42);
	s_in2(9,42)            <= s_out2(10,43);
	s_locks_lower_in(9,42) <= s_locks_lower_out(10,42);

		normal_cell_9_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,43),
			fetch              => s_fetch(9,43),
			data_in            => s_data_in(9,43),
			data_out           => s_data_out(9,43),
			out1               => s_out1(9,43),
			out2               => s_out2(9,43),
			lock_lower_row_out => s_locks_lower_out(9,43),
			lock_lower_row_in  => s_locks_lower_in(9,43),
			in1                => s_in1(9,43),
			in2                => s_in2(9,43),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(43)
		);
	s_in1(9,43)            <= s_out1(10,43);
	s_in2(9,43)            <= s_out2(10,44);
	s_locks_lower_in(9,43) <= s_locks_lower_out(10,43);

		normal_cell_9_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,44),
			fetch              => s_fetch(9,44),
			data_in            => s_data_in(9,44),
			data_out           => s_data_out(9,44),
			out1               => s_out1(9,44),
			out2               => s_out2(9,44),
			lock_lower_row_out => s_locks_lower_out(9,44),
			lock_lower_row_in  => s_locks_lower_in(9,44),
			in1                => s_in1(9,44),
			in2                => s_in2(9,44),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(44)
		);
	s_in1(9,44)            <= s_out1(10,44);
	s_in2(9,44)            <= s_out2(10,45);
	s_locks_lower_in(9,44) <= s_locks_lower_out(10,44);

		normal_cell_9_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,45),
			fetch              => s_fetch(9,45),
			data_in            => s_data_in(9,45),
			data_out           => s_data_out(9,45),
			out1               => s_out1(9,45),
			out2               => s_out2(9,45),
			lock_lower_row_out => s_locks_lower_out(9,45),
			lock_lower_row_in  => s_locks_lower_in(9,45),
			in1                => s_in1(9,45),
			in2                => s_in2(9,45),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(45)
		);
	s_in1(9,45)            <= s_out1(10,45);
	s_in2(9,45)            <= s_out2(10,46);
	s_locks_lower_in(9,45) <= s_locks_lower_out(10,45);

		normal_cell_9_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,46),
			fetch              => s_fetch(9,46),
			data_in            => s_data_in(9,46),
			data_out           => s_data_out(9,46),
			out1               => s_out1(9,46),
			out2               => s_out2(9,46),
			lock_lower_row_out => s_locks_lower_out(9,46),
			lock_lower_row_in  => s_locks_lower_in(9,46),
			in1                => s_in1(9,46),
			in2                => s_in2(9,46),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(46)
		);
	s_in1(9,46)            <= s_out1(10,46);
	s_in2(9,46)            <= s_out2(10,47);
	s_locks_lower_in(9,46) <= s_locks_lower_out(10,46);

		normal_cell_9_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,47),
			fetch              => s_fetch(9,47),
			data_in            => s_data_in(9,47),
			data_out           => s_data_out(9,47),
			out1               => s_out1(9,47),
			out2               => s_out2(9,47),
			lock_lower_row_out => s_locks_lower_out(9,47),
			lock_lower_row_in  => s_locks_lower_in(9,47),
			in1                => s_in1(9,47),
			in2                => s_in2(9,47),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(47)
		);
	s_in1(9,47)            <= s_out1(10,47);
	s_in2(9,47)            <= s_out2(10,48);
	s_locks_lower_in(9,47) <= s_locks_lower_out(10,47);

		normal_cell_9_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,48),
			fetch              => s_fetch(9,48),
			data_in            => s_data_in(9,48),
			data_out           => s_data_out(9,48),
			out1               => s_out1(9,48),
			out2               => s_out2(9,48),
			lock_lower_row_out => s_locks_lower_out(9,48),
			lock_lower_row_in  => s_locks_lower_in(9,48),
			in1                => s_in1(9,48),
			in2                => s_in2(9,48),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(48)
		);
	s_in1(9,48)            <= s_out1(10,48);
	s_in2(9,48)            <= s_out2(10,49);
	s_locks_lower_in(9,48) <= s_locks_lower_out(10,48);

		normal_cell_9_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,49),
			fetch              => s_fetch(9,49),
			data_in            => s_data_in(9,49),
			data_out           => s_data_out(9,49),
			out1               => s_out1(9,49),
			out2               => s_out2(9,49),
			lock_lower_row_out => s_locks_lower_out(9,49),
			lock_lower_row_in  => s_locks_lower_in(9,49),
			in1                => s_in1(9,49),
			in2                => s_in2(9,49),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(49)
		);
	s_in1(9,49)            <= s_out1(10,49);
	s_in2(9,49)            <= s_out2(10,50);
	s_locks_lower_in(9,49) <= s_locks_lower_out(10,49);

		normal_cell_9_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,50),
			fetch              => s_fetch(9,50),
			data_in            => s_data_in(9,50),
			data_out           => s_data_out(9,50),
			out1               => s_out1(9,50),
			out2               => s_out2(9,50),
			lock_lower_row_out => s_locks_lower_out(9,50),
			lock_lower_row_in  => s_locks_lower_in(9,50),
			in1                => s_in1(9,50),
			in2                => s_in2(9,50),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(50)
		);
	s_in1(9,50)            <= s_out1(10,50);
	s_in2(9,50)            <= s_out2(10,51);
	s_locks_lower_in(9,50) <= s_locks_lower_out(10,50);

		normal_cell_9_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,51),
			fetch              => s_fetch(9,51),
			data_in            => s_data_in(9,51),
			data_out           => s_data_out(9,51),
			out1               => s_out1(9,51),
			out2               => s_out2(9,51),
			lock_lower_row_out => s_locks_lower_out(9,51),
			lock_lower_row_in  => s_locks_lower_in(9,51),
			in1                => s_in1(9,51),
			in2                => s_in2(9,51),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(51)
		);
	s_in1(9,51)            <= s_out1(10,51);
	s_in2(9,51)            <= s_out2(10,52);
	s_locks_lower_in(9,51) <= s_locks_lower_out(10,51);

		normal_cell_9_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,52),
			fetch              => s_fetch(9,52),
			data_in            => s_data_in(9,52),
			data_out           => s_data_out(9,52),
			out1               => s_out1(9,52),
			out2               => s_out2(9,52),
			lock_lower_row_out => s_locks_lower_out(9,52),
			lock_lower_row_in  => s_locks_lower_in(9,52),
			in1                => s_in1(9,52),
			in2                => s_in2(9,52),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(52)
		);
	s_in1(9,52)            <= s_out1(10,52);
	s_in2(9,52)            <= s_out2(10,53);
	s_locks_lower_in(9,52) <= s_locks_lower_out(10,52);

		normal_cell_9_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,53),
			fetch              => s_fetch(9,53),
			data_in            => s_data_in(9,53),
			data_out           => s_data_out(9,53),
			out1               => s_out1(9,53),
			out2               => s_out2(9,53),
			lock_lower_row_out => s_locks_lower_out(9,53),
			lock_lower_row_in  => s_locks_lower_in(9,53),
			in1                => s_in1(9,53),
			in2                => s_in2(9,53),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(53)
		);
	s_in1(9,53)            <= s_out1(10,53);
	s_in2(9,53)            <= s_out2(10,54);
	s_locks_lower_in(9,53) <= s_locks_lower_out(10,53);

		normal_cell_9_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,54),
			fetch              => s_fetch(9,54),
			data_in            => s_data_in(9,54),
			data_out           => s_data_out(9,54),
			out1               => s_out1(9,54),
			out2               => s_out2(9,54),
			lock_lower_row_out => s_locks_lower_out(9,54),
			lock_lower_row_in  => s_locks_lower_in(9,54),
			in1                => s_in1(9,54),
			in2                => s_in2(9,54),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(54)
		);
	s_in1(9,54)            <= s_out1(10,54);
	s_in2(9,54)            <= s_out2(10,55);
	s_locks_lower_in(9,54) <= s_locks_lower_out(10,54);

		normal_cell_9_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,55),
			fetch              => s_fetch(9,55),
			data_in            => s_data_in(9,55),
			data_out           => s_data_out(9,55),
			out1               => s_out1(9,55),
			out2               => s_out2(9,55),
			lock_lower_row_out => s_locks_lower_out(9,55),
			lock_lower_row_in  => s_locks_lower_in(9,55),
			in1                => s_in1(9,55),
			in2                => s_in2(9,55),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(55)
		);
	s_in1(9,55)            <= s_out1(10,55);
	s_in2(9,55)            <= s_out2(10,56);
	s_locks_lower_in(9,55) <= s_locks_lower_out(10,55);

		normal_cell_9_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,56),
			fetch              => s_fetch(9,56),
			data_in            => s_data_in(9,56),
			data_out           => s_data_out(9,56),
			out1               => s_out1(9,56),
			out2               => s_out2(9,56),
			lock_lower_row_out => s_locks_lower_out(9,56),
			lock_lower_row_in  => s_locks_lower_in(9,56),
			in1                => s_in1(9,56),
			in2                => s_in2(9,56),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(56)
		);
	s_in1(9,56)            <= s_out1(10,56);
	s_in2(9,56)            <= s_out2(10,57);
	s_locks_lower_in(9,56) <= s_locks_lower_out(10,56);

		normal_cell_9_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,57),
			fetch              => s_fetch(9,57),
			data_in            => s_data_in(9,57),
			data_out           => s_data_out(9,57),
			out1               => s_out1(9,57),
			out2               => s_out2(9,57),
			lock_lower_row_out => s_locks_lower_out(9,57),
			lock_lower_row_in  => s_locks_lower_in(9,57),
			in1                => s_in1(9,57),
			in2                => s_in2(9,57),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(57)
		);
	s_in1(9,57)            <= s_out1(10,57);
	s_in2(9,57)            <= s_out2(10,58);
	s_locks_lower_in(9,57) <= s_locks_lower_out(10,57);

		normal_cell_9_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,58),
			fetch              => s_fetch(9,58),
			data_in            => s_data_in(9,58),
			data_out           => s_data_out(9,58),
			out1               => s_out1(9,58),
			out2               => s_out2(9,58),
			lock_lower_row_out => s_locks_lower_out(9,58),
			lock_lower_row_in  => s_locks_lower_in(9,58),
			in1                => s_in1(9,58),
			in2                => s_in2(9,58),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(58)
		);
	s_in1(9,58)            <= s_out1(10,58);
	s_in2(9,58)            <= s_out2(10,59);
	s_locks_lower_in(9,58) <= s_locks_lower_out(10,58);

		normal_cell_9_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,59),
			fetch              => s_fetch(9,59),
			data_in            => s_data_in(9,59),
			data_out           => s_data_out(9,59),
			out1               => s_out1(9,59),
			out2               => s_out2(9,59),
			lock_lower_row_out => s_locks_lower_out(9,59),
			lock_lower_row_in  => s_locks_lower_in(9,59),
			in1                => s_in1(9,59),
			in2                => s_in2(9,59),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(59)
		);
	s_in1(9,59)            <= s_out1(10,59);
	s_in2(9,59)            <= s_out2(10,60);
	s_locks_lower_in(9,59) <= s_locks_lower_out(10,59);

		last_col_cell_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(9,60),
			fetch              => s_fetch(9,60),
			data_in            => s_data_in(9,60),
			data_out           => s_data_out(9,60),
			out1               => s_out1(9,60),
			out2               => s_out2(9,60),
			lock_lower_row_out => s_locks_lower_out(9,60),
			lock_lower_row_in  => s_locks_lower_in(9,60),
			in1                => s_in1(9,60),
			in2                => (others => '0'),
			lock_row           => s_locks(9),
			piv_found          => s_piv_found,
			row_data           => s_row_data(9),
			col_data           => s_col_data(60)
		);
	s_in1(9,60)            <= s_out1(10,60);
	s_locks_lower_in(9,60) <= s_locks_lower_out(10,60);

		normal_cell_10_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,1),
			fetch              => s_fetch(10,1),
			data_in            => s_data_in(10,1),
			data_out           => s_data_out(10,1),
			out1               => s_out1(10,1),
			out2               => s_out2(10,1),
			lock_lower_row_out => s_locks_lower_out(10,1),
			lock_lower_row_in  => s_locks_lower_in(10,1),
			in1                => s_in1(10,1),
			in2                => s_in2(10,1),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(1)
		);
	s_in1(10,1)            <= s_out1(11,1);
	s_in2(10,1)            <= s_out2(11,2);
	s_locks_lower_in(10,1) <= s_locks_lower_out(11,1);

		normal_cell_10_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,2),
			fetch              => s_fetch(10,2),
			data_in            => s_data_in(10,2),
			data_out           => s_data_out(10,2),
			out1               => s_out1(10,2),
			out2               => s_out2(10,2),
			lock_lower_row_out => s_locks_lower_out(10,2),
			lock_lower_row_in  => s_locks_lower_in(10,2),
			in1                => s_in1(10,2),
			in2                => s_in2(10,2),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(2)
		);
	s_in1(10,2)            <= s_out1(11,2);
	s_in2(10,2)            <= s_out2(11,3);
	s_locks_lower_in(10,2) <= s_locks_lower_out(11,2);

		normal_cell_10_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,3),
			fetch              => s_fetch(10,3),
			data_in            => s_data_in(10,3),
			data_out           => s_data_out(10,3),
			out1               => s_out1(10,3),
			out2               => s_out2(10,3),
			lock_lower_row_out => s_locks_lower_out(10,3),
			lock_lower_row_in  => s_locks_lower_in(10,3),
			in1                => s_in1(10,3),
			in2                => s_in2(10,3),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(3)
		);
	s_in1(10,3)            <= s_out1(11,3);
	s_in2(10,3)            <= s_out2(11,4);
	s_locks_lower_in(10,3) <= s_locks_lower_out(11,3);

		normal_cell_10_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,4),
			fetch              => s_fetch(10,4),
			data_in            => s_data_in(10,4),
			data_out           => s_data_out(10,4),
			out1               => s_out1(10,4),
			out2               => s_out2(10,4),
			lock_lower_row_out => s_locks_lower_out(10,4),
			lock_lower_row_in  => s_locks_lower_in(10,4),
			in1                => s_in1(10,4),
			in2                => s_in2(10,4),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(4)
		);
	s_in1(10,4)            <= s_out1(11,4);
	s_in2(10,4)            <= s_out2(11,5);
	s_locks_lower_in(10,4) <= s_locks_lower_out(11,4);

		normal_cell_10_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,5),
			fetch              => s_fetch(10,5),
			data_in            => s_data_in(10,5),
			data_out           => s_data_out(10,5),
			out1               => s_out1(10,5),
			out2               => s_out2(10,5),
			lock_lower_row_out => s_locks_lower_out(10,5),
			lock_lower_row_in  => s_locks_lower_in(10,5),
			in1                => s_in1(10,5),
			in2                => s_in2(10,5),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(5)
		);
	s_in1(10,5)            <= s_out1(11,5);
	s_in2(10,5)            <= s_out2(11,6);
	s_locks_lower_in(10,5) <= s_locks_lower_out(11,5);

		normal_cell_10_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,6),
			fetch              => s_fetch(10,6),
			data_in            => s_data_in(10,6),
			data_out           => s_data_out(10,6),
			out1               => s_out1(10,6),
			out2               => s_out2(10,6),
			lock_lower_row_out => s_locks_lower_out(10,6),
			lock_lower_row_in  => s_locks_lower_in(10,6),
			in1                => s_in1(10,6),
			in2                => s_in2(10,6),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(6)
		);
	s_in1(10,6)            <= s_out1(11,6);
	s_in2(10,6)            <= s_out2(11,7);
	s_locks_lower_in(10,6) <= s_locks_lower_out(11,6);

		normal_cell_10_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,7),
			fetch              => s_fetch(10,7),
			data_in            => s_data_in(10,7),
			data_out           => s_data_out(10,7),
			out1               => s_out1(10,7),
			out2               => s_out2(10,7),
			lock_lower_row_out => s_locks_lower_out(10,7),
			lock_lower_row_in  => s_locks_lower_in(10,7),
			in1                => s_in1(10,7),
			in2                => s_in2(10,7),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(7)
		);
	s_in1(10,7)            <= s_out1(11,7);
	s_in2(10,7)            <= s_out2(11,8);
	s_locks_lower_in(10,7) <= s_locks_lower_out(11,7);

		normal_cell_10_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,8),
			fetch              => s_fetch(10,8),
			data_in            => s_data_in(10,8),
			data_out           => s_data_out(10,8),
			out1               => s_out1(10,8),
			out2               => s_out2(10,8),
			lock_lower_row_out => s_locks_lower_out(10,8),
			lock_lower_row_in  => s_locks_lower_in(10,8),
			in1                => s_in1(10,8),
			in2                => s_in2(10,8),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(8)
		);
	s_in1(10,8)            <= s_out1(11,8);
	s_in2(10,8)            <= s_out2(11,9);
	s_locks_lower_in(10,8) <= s_locks_lower_out(11,8);

		normal_cell_10_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,9),
			fetch              => s_fetch(10,9),
			data_in            => s_data_in(10,9),
			data_out           => s_data_out(10,9),
			out1               => s_out1(10,9),
			out2               => s_out2(10,9),
			lock_lower_row_out => s_locks_lower_out(10,9),
			lock_lower_row_in  => s_locks_lower_in(10,9),
			in1                => s_in1(10,9),
			in2                => s_in2(10,9),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(9)
		);
	s_in1(10,9)            <= s_out1(11,9);
	s_in2(10,9)            <= s_out2(11,10);
	s_locks_lower_in(10,9) <= s_locks_lower_out(11,9);

		normal_cell_10_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,10),
			fetch              => s_fetch(10,10),
			data_in            => s_data_in(10,10),
			data_out           => s_data_out(10,10),
			out1               => s_out1(10,10),
			out2               => s_out2(10,10),
			lock_lower_row_out => s_locks_lower_out(10,10),
			lock_lower_row_in  => s_locks_lower_in(10,10),
			in1                => s_in1(10,10),
			in2                => s_in2(10,10),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(10)
		);
	s_in1(10,10)            <= s_out1(11,10);
	s_in2(10,10)            <= s_out2(11,11);
	s_locks_lower_in(10,10) <= s_locks_lower_out(11,10);

		normal_cell_10_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,11),
			fetch              => s_fetch(10,11),
			data_in            => s_data_in(10,11),
			data_out           => s_data_out(10,11),
			out1               => s_out1(10,11),
			out2               => s_out2(10,11),
			lock_lower_row_out => s_locks_lower_out(10,11),
			lock_lower_row_in  => s_locks_lower_in(10,11),
			in1                => s_in1(10,11),
			in2                => s_in2(10,11),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(11)
		);
	s_in1(10,11)            <= s_out1(11,11);
	s_in2(10,11)            <= s_out2(11,12);
	s_locks_lower_in(10,11) <= s_locks_lower_out(11,11);

		normal_cell_10_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,12),
			fetch              => s_fetch(10,12),
			data_in            => s_data_in(10,12),
			data_out           => s_data_out(10,12),
			out1               => s_out1(10,12),
			out2               => s_out2(10,12),
			lock_lower_row_out => s_locks_lower_out(10,12),
			lock_lower_row_in  => s_locks_lower_in(10,12),
			in1                => s_in1(10,12),
			in2                => s_in2(10,12),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(12)
		);
	s_in1(10,12)            <= s_out1(11,12);
	s_in2(10,12)            <= s_out2(11,13);
	s_locks_lower_in(10,12) <= s_locks_lower_out(11,12);

		normal_cell_10_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,13),
			fetch              => s_fetch(10,13),
			data_in            => s_data_in(10,13),
			data_out           => s_data_out(10,13),
			out1               => s_out1(10,13),
			out2               => s_out2(10,13),
			lock_lower_row_out => s_locks_lower_out(10,13),
			lock_lower_row_in  => s_locks_lower_in(10,13),
			in1                => s_in1(10,13),
			in2                => s_in2(10,13),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(13)
		);
	s_in1(10,13)            <= s_out1(11,13);
	s_in2(10,13)            <= s_out2(11,14);
	s_locks_lower_in(10,13) <= s_locks_lower_out(11,13);

		normal_cell_10_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,14),
			fetch              => s_fetch(10,14),
			data_in            => s_data_in(10,14),
			data_out           => s_data_out(10,14),
			out1               => s_out1(10,14),
			out2               => s_out2(10,14),
			lock_lower_row_out => s_locks_lower_out(10,14),
			lock_lower_row_in  => s_locks_lower_in(10,14),
			in1                => s_in1(10,14),
			in2                => s_in2(10,14),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(14)
		);
	s_in1(10,14)            <= s_out1(11,14);
	s_in2(10,14)            <= s_out2(11,15);
	s_locks_lower_in(10,14) <= s_locks_lower_out(11,14);

		normal_cell_10_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,15),
			fetch              => s_fetch(10,15),
			data_in            => s_data_in(10,15),
			data_out           => s_data_out(10,15),
			out1               => s_out1(10,15),
			out2               => s_out2(10,15),
			lock_lower_row_out => s_locks_lower_out(10,15),
			lock_lower_row_in  => s_locks_lower_in(10,15),
			in1                => s_in1(10,15),
			in2                => s_in2(10,15),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(15)
		);
	s_in1(10,15)            <= s_out1(11,15);
	s_in2(10,15)            <= s_out2(11,16);
	s_locks_lower_in(10,15) <= s_locks_lower_out(11,15);

		normal_cell_10_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,16),
			fetch              => s_fetch(10,16),
			data_in            => s_data_in(10,16),
			data_out           => s_data_out(10,16),
			out1               => s_out1(10,16),
			out2               => s_out2(10,16),
			lock_lower_row_out => s_locks_lower_out(10,16),
			lock_lower_row_in  => s_locks_lower_in(10,16),
			in1                => s_in1(10,16),
			in2                => s_in2(10,16),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(16)
		);
	s_in1(10,16)            <= s_out1(11,16);
	s_in2(10,16)            <= s_out2(11,17);
	s_locks_lower_in(10,16) <= s_locks_lower_out(11,16);

		normal_cell_10_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,17),
			fetch              => s_fetch(10,17),
			data_in            => s_data_in(10,17),
			data_out           => s_data_out(10,17),
			out1               => s_out1(10,17),
			out2               => s_out2(10,17),
			lock_lower_row_out => s_locks_lower_out(10,17),
			lock_lower_row_in  => s_locks_lower_in(10,17),
			in1                => s_in1(10,17),
			in2                => s_in2(10,17),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(17)
		);
	s_in1(10,17)            <= s_out1(11,17);
	s_in2(10,17)            <= s_out2(11,18);
	s_locks_lower_in(10,17) <= s_locks_lower_out(11,17);

		normal_cell_10_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,18),
			fetch              => s_fetch(10,18),
			data_in            => s_data_in(10,18),
			data_out           => s_data_out(10,18),
			out1               => s_out1(10,18),
			out2               => s_out2(10,18),
			lock_lower_row_out => s_locks_lower_out(10,18),
			lock_lower_row_in  => s_locks_lower_in(10,18),
			in1                => s_in1(10,18),
			in2                => s_in2(10,18),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(18)
		);
	s_in1(10,18)            <= s_out1(11,18);
	s_in2(10,18)            <= s_out2(11,19);
	s_locks_lower_in(10,18) <= s_locks_lower_out(11,18);

		normal_cell_10_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,19),
			fetch              => s_fetch(10,19),
			data_in            => s_data_in(10,19),
			data_out           => s_data_out(10,19),
			out1               => s_out1(10,19),
			out2               => s_out2(10,19),
			lock_lower_row_out => s_locks_lower_out(10,19),
			lock_lower_row_in  => s_locks_lower_in(10,19),
			in1                => s_in1(10,19),
			in2                => s_in2(10,19),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(19)
		);
	s_in1(10,19)            <= s_out1(11,19);
	s_in2(10,19)            <= s_out2(11,20);
	s_locks_lower_in(10,19) <= s_locks_lower_out(11,19);

		normal_cell_10_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,20),
			fetch              => s_fetch(10,20),
			data_in            => s_data_in(10,20),
			data_out           => s_data_out(10,20),
			out1               => s_out1(10,20),
			out2               => s_out2(10,20),
			lock_lower_row_out => s_locks_lower_out(10,20),
			lock_lower_row_in  => s_locks_lower_in(10,20),
			in1                => s_in1(10,20),
			in2                => s_in2(10,20),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(20)
		);
	s_in1(10,20)            <= s_out1(11,20);
	s_in2(10,20)            <= s_out2(11,21);
	s_locks_lower_in(10,20) <= s_locks_lower_out(11,20);

		normal_cell_10_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,21),
			fetch              => s_fetch(10,21),
			data_in            => s_data_in(10,21),
			data_out           => s_data_out(10,21),
			out1               => s_out1(10,21),
			out2               => s_out2(10,21),
			lock_lower_row_out => s_locks_lower_out(10,21),
			lock_lower_row_in  => s_locks_lower_in(10,21),
			in1                => s_in1(10,21),
			in2                => s_in2(10,21),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(21)
		);
	s_in1(10,21)            <= s_out1(11,21);
	s_in2(10,21)            <= s_out2(11,22);
	s_locks_lower_in(10,21) <= s_locks_lower_out(11,21);

		normal_cell_10_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,22),
			fetch              => s_fetch(10,22),
			data_in            => s_data_in(10,22),
			data_out           => s_data_out(10,22),
			out1               => s_out1(10,22),
			out2               => s_out2(10,22),
			lock_lower_row_out => s_locks_lower_out(10,22),
			lock_lower_row_in  => s_locks_lower_in(10,22),
			in1                => s_in1(10,22),
			in2                => s_in2(10,22),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(22)
		);
	s_in1(10,22)            <= s_out1(11,22);
	s_in2(10,22)            <= s_out2(11,23);
	s_locks_lower_in(10,22) <= s_locks_lower_out(11,22);

		normal_cell_10_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,23),
			fetch              => s_fetch(10,23),
			data_in            => s_data_in(10,23),
			data_out           => s_data_out(10,23),
			out1               => s_out1(10,23),
			out2               => s_out2(10,23),
			lock_lower_row_out => s_locks_lower_out(10,23),
			lock_lower_row_in  => s_locks_lower_in(10,23),
			in1                => s_in1(10,23),
			in2                => s_in2(10,23),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(23)
		);
	s_in1(10,23)            <= s_out1(11,23);
	s_in2(10,23)            <= s_out2(11,24);
	s_locks_lower_in(10,23) <= s_locks_lower_out(11,23);

		normal_cell_10_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,24),
			fetch              => s_fetch(10,24),
			data_in            => s_data_in(10,24),
			data_out           => s_data_out(10,24),
			out1               => s_out1(10,24),
			out2               => s_out2(10,24),
			lock_lower_row_out => s_locks_lower_out(10,24),
			lock_lower_row_in  => s_locks_lower_in(10,24),
			in1                => s_in1(10,24),
			in2                => s_in2(10,24),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(24)
		);
	s_in1(10,24)            <= s_out1(11,24);
	s_in2(10,24)            <= s_out2(11,25);
	s_locks_lower_in(10,24) <= s_locks_lower_out(11,24);

		normal_cell_10_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,25),
			fetch              => s_fetch(10,25),
			data_in            => s_data_in(10,25),
			data_out           => s_data_out(10,25),
			out1               => s_out1(10,25),
			out2               => s_out2(10,25),
			lock_lower_row_out => s_locks_lower_out(10,25),
			lock_lower_row_in  => s_locks_lower_in(10,25),
			in1                => s_in1(10,25),
			in2                => s_in2(10,25),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(25)
		);
	s_in1(10,25)            <= s_out1(11,25);
	s_in2(10,25)            <= s_out2(11,26);
	s_locks_lower_in(10,25) <= s_locks_lower_out(11,25);

		normal_cell_10_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,26),
			fetch              => s_fetch(10,26),
			data_in            => s_data_in(10,26),
			data_out           => s_data_out(10,26),
			out1               => s_out1(10,26),
			out2               => s_out2(10,26),
			lock_lower_row_out => s_locks_lower_out(10,26),
			lock_lower_row_in  => s_locks_lower_in(10,26),
			in1                => s_in1(10,26),
			in2                => s_in2(10,26),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(26)
		);
	s_in1(10,26)            <= s_out1(11,26);
	s_in2(10,26)            <= s_out2(11,27);
	s_locks_lower_in(10,26) <= s_locks_lower_out(11,26);

		normal_cell_10_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,27),
			fetch              => s_fetch(10,27),
			data_in            => s_data_in(10,27),
			data_out           => s_data_out(10,27),
			out1               => s_out1(10,27),
			out2               => s_out2(10,27),
			lock_lower_row_out => s_locks_lower_out(10,27),
			lock_lower_row_in  => s_locks_lower_in(10,27),
			in1                => s_in1(10,27),
			in2                => s_in2(10,27),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(27)
		);
	s_in1(10,27)            <= s_out1(11,27);
	s_in2(10,27)            <= s_out2(11,28);
	s_locks_lower_in(10,27) <= s_locks_lower_out(11,27);

		normal_cell_10_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,28),
			fetch              => s_fetch(10,28),
			data_in            => s_data_in(10,28),
			data_out           => s_data_out(10,28),
			out1               => s_out1(10,28),
			out2               => s_out2(10,28),
			lock_lower_row_out => s_locks_lower_out(10,28),
			lock_lower_row_in  => s_locks_lower_in(10,28),
			in1                => s_in1(10,28),
			in2                => s_in2(10,28),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(28)
		);
	s_in1(10,28)            <= s_out1(11,28);
	s_in2(10,28)            <= s_out2(11,29);
	s_locks_lower_in(10,28) <= s_locks_lower_out(11,28);

		normal_cell_10_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,29),
			fetch              => s_fetch(10,29),
			data_in            => s_data_in(10,29),
			data_out           => s_data_out(10,29),
			out1               => s_out1(10,29),
			out2               => s_out2(10,29),
			lock_lower_row_out => s_locks_lower_out(10,29),
			lock_lower_row_in  => s_locks_lower_in(10,29),
			in1                => s_in1(10,29),
			in2                => s_in2(10,29),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(29)
		);
	s_in1(10,29)            <= s_out1(11,29);
	s_in2(10,29)            <= s_out2(11,30);
	s_locks_lower_in(10,29) <= s_locks_lower_out(11,29);

		normal_cell_10_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,30),
			fetch              => s_fetch(10,30),
			data_in            => s_data_in(10,30),
			data_out           => s_data_out(10,30),
			out1               => s_out1(10,30),
			out2               => s_out2(10,30),
			lock_lower_row_out => s_locks_lower_out(10,30),
			lock_lower_row_in  => s_locks_lower_in(10,30),
			in1                => s_in1(10,30),
			in2                => s_in2(10,30),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(30)
		);
	s_in1(10,30)            <= s_out1(11,30);
	s_in2(10,30)            <= s_out2(11,31);
	s_locks_lower_in(10,30) <= s_locks_lower_out(11,30);

		normal_cell_10_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,31),
			fetch              => s_fetch(10,31),
			data_in            => s_data_in(10,31),
			data_out           => s_data_out(10,31),
			out1               => s_out1(10,31),
			out2               => s_out2(10,31),
			lock_lower_row_out => s_locks_lower_out(10,31),
			lock_lower_row_in  => s_locks_lower_in(10,31),
			in1                => s_in1(10,31),
			in2                => s_in2(10,31),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(31)
		);
	s_in1(10,31)            <= s_out1(11,31);
	s_in2(10,31)            <= s_out2(11,32);
	s_locks_lower_in(10,31) <= s_locks_lower_out(11,31);

		normal_cell_10_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,32),
			fetch              => s_fetch(10,32),
			data_in            => s_data_in(10,32),
			data_out           => s_data_out(10,32),
			out1               => s_out1(10,32),
			out2               => s_out2(10,32),
			lock_lower_row_out => s_locks_lower_out(10,32),
			lock_lower_row_in  => s_locks_lower_in(10,32),
			in1                => s_in1(10,32),
			in2                => s_in2(10,32),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(32)
		);
	s_in1(10,32)            <= s_out1(11,32);
	s_in2(10,32)            <= s_out2(11,33);
	s_locks_lower_in(10,32) <= s_locks_lower_out(11,32);

		normal_cell_10_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,33),
			fetch              => s_fetch(10,33),
			data_in            => s_data_in(10,33),
			data_out           => s_data_out(10,33),
			out1               => s_out1(10,33),
			out2               => s_out2(10,33),
			lock_lower_row_out => s_locks_lower_out(10,33),
			lock_lower_row_in  => s_locks_lower_in(10,33),
			in1                => s_in1(10,33),
			in2                => s_in2(10,33),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(33)
		);
	s_in1(10,33)            <= s_out1(11,33);
	s_in2(10,33)            <= s_out2(11,34);
	s_locks_lower_in(10,33) <= s_locks_lower_out(11,33);

		normal_cell_10_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,34),
			fetch              => s_fetch(10,34),
			data_in            => s_data_in(10,34),
			data_out           => s_data_out(10,34),
			out1               => s_out1(10,34),
			out2               => s_out2(10,34),
			lock_lower_row_out => s_locks_lower_out(10,34),
			lock_lower_row_in  => s_locks_lower_in(10,34),
			in1                => s_in1(10,34),
			in2                => s_in2(10,34),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(34)
		);
	s_in1(10,34)            <= s_out1(11,34);
	s_in2(10,34)            <= s_out2(11,35);
	s_locks_lower_in(10,34) <= s_locks_lower_out(11,34);

		normal_cell_10_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,35),
			fetch              => s_fetch(10,35),
			data_in            => s_data_in(10,35),
			data_out           => s_data_out(10,35),
			out1               => s_out1(10,35),
			out2               => s_out2(10,35),
			lock_lower_row_out => s_locks_lower_out(10,35),
			lock_lower_row_in  => s_locks_lower_in(10,35),
			in1                => s_in1(10,35),
			in2                => s_in2(10,35),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(35)
		);
	s_in1(10,35)            <= s_out1(11,35);
	s_in2(10,35)            <= s_out2(11,36);
	s_locks_lower_in(10,35) <= s_locks_lower_out(11,35);

		normal_cell_10_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,36),
			fetch              => s_fetch(10,36),
			data_in            => s_data_in(10,36),
			data_out           => s_data_out(10,36),
			out1               => s_out1(10,36),
			out2               => s_out2(10,36),
			lock_lower_row_out => s_locks_lower_out(10,36),
			lock_lower_row_in  => s_locks_lower_in(10,36),
			in1                => s_in1(10,36),
			in2                => s_in2(10,36),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(36)
		);
	s_in1(10,36)            <= s_out1(11,36);
	s_in2(10,36)            <= s_out2(11,37);
	s_locks_lower_in(10,36) <= s_locks_lower_out(11,36);

		normal_cell_10_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,37),
			fetch              => s_fetch(10,37),
			data_in            => s_data_in(10,37),
			data_out           => s_data_out(10,37),
			out1               => s_out1(10,37),
			out2               => s_out2(10,37),
			lock_lower_row_out => s_locks_lower_out(10,37),
			lock_lower_row_in  => s_locks_lower_in(10,37),
			in1                => s_in1(10,37),
			in2                => s_in2(10,37),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(37)
		);
	s_in1(10,37)            <= s_out1(11,37);
	s_in2(10,37)            <= s_out2(11,38);
	s_locks_lower_in(10,37) <= s_locks_lower_out(11,37);

		normal_cell_10_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,38),
			fetch              => s_fetch(10,38),
			data_in            => s_data_in(10,38),
			data_out           => s_data_out(10,38),
			out1               => s_out1(10,38),
			out2               => s_out2(10,38),
			lock_lower_row_out => s_locks_lower_out(10,38),
			lock_lower_row_in  => s_locks_lower_in(10,38),
			in1                => s_in1(10,38),
			in2                => s_in2(10,38),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(38)
		);
	s_in1(10,38)            <= s_out1(11,38);
	s_in2(10,38)            <= s_out2(11,39);
	s_locks_lower_in(10,38) <= s_locks_lower_out(11,38);

		normal_cell_10_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,39),
			fetch              => s_fetch(10,39),
			data_in            => s_data_in(10,39),
			data_out           => s_data_out(10,39),
			out1               => s_out1(10,39),
			out2               => s_out2(10,39),
			lock_lower_row_out => s_locks_lower_out(10,39),
			lock_lower_row_in  => s_locks_lower_in(10,39),
			in1                => s_in1(10,39),
			in2                => s_in2(10,39),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(39)
		);
	s_in1(10,39)            <= s_out1(11,39);
	s_in2(10,39)            <= s_out2(11,40);
	s_locks_lower_in(10,39) <= s_locks_lower_out(11,39);

		normal_cell_10_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,40),
			fetch              => s_fetch(10,40),
			data_in            => s_data_in(10,40),
			data_out           => s_data_out(10,40),
			out1               => s_out1(10,40),
			out2               => s_out2(10,40),
			lock_lower_row_out => s_locks_lower_out(10,40),
			lock_lower_row_in  => s_locks_lower_in(10,40),
			in1                => s_in1(10,40),
			in2                => s_in2(10,40),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(40)
		);
	s_in1(10,40)            <= s_out1(11,40);
	s_in2(10,40)            <= s_out2(11,41);
	s_locks_lower_in(10,40) <= s_locks_lower_out(11,40);

		normal_cell_10_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,41),
			fetch              => s_fetch(10,41),
			data_in            => s_data_in(10,41),
			data_out           => s_data_out(10,41),
			out1               => s_out1(10,41),
			out2               => s_out2(10,41),
			lock_lower_row_out => s_locks_lower_out(10,41),
			lock_lower_row_in  => s_locks_lower_in(10,41),
			in1                => s_in1(10,41),
			in2                => s_in2(10,41),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(41)
		);
	s_in1(10,41)            <= s_out1(11,41);
	s_in2(10,41)            <= s_out2(11,42);
	s_locks_lower_in(10,41) <= s_locks_lower_out(11,41);

		normal_cell_10_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,42),
			fetch              => s_fetch(10,42),
			data_in            => s_data_in(10,42),
			data_out           => s_data_out(10,42),
			out1               => s_out1(10,42),
			out2               => s_out2(10,42),
			lock_lower_row_out => s_locks_lower_out(10,42),
			lock_lower_row_in  => s_locks_lower_in(10,42),
			in1                => s_in1(10,42),
			in2                => s_in2(10,42),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(42)
		);
	s_in1(10,42)            <= s_out1(11,42);
	s_in2(10,42)            <= s_out2(11,43);
	s_locks_lower_in(10,42) <= s_locks_lower_out(11,42);

		normal_cell_10_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,43),
			fetch              => s_fetch(10,43),
			data_in            => s_data_in(10,43),
			data_out           => s_data_out(10,43),
			out1               => s_out1(10,43),
			out2               => s_out2(10,43),
			lock_lower_row_out => s_locks_lower_out(10,43),
			lock_lower_row_in  => s_locks_lower_in(10,43),
			in1                => s_in1(10,43),
			in2                => s_in2(10,43),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(43)
		);
	s_in1(10,43)            <= s_out1(11,43);
	s_in2(10,43)            <= s_out2(11,44);
	s_locks_lower_in(10,43) <= s_locks_lower_out(11,43);

		normal_cell_10_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,44),
			fetch              => s_fetch(10,44),
			data_in            => s_data_in(10,44),
			data_out           => s_data_out(10,44),
			out1               => s_out1(10,44),
			out2               => s_out2(10,44),
			lock_lower_row_out => s_locks_lower_out(10,44),
			lock_lower_row_in  => s_locks_lower_in(10,44),
			in1                => s_in1(10,44),
			in2                => s_in2(10,44),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(44)
		);
	s_in1(10,44)            <= s_out1(11,44);
	s_in2(10,44)            <= s_out2(11,45);
	s_locks_lower_in(10,44) <= s_locks_lower_out(11,44);

		normal_cell_10_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,45),
			fetch              => s_fetch(10,45),
			data_in            => s_data_in(10,45),
			data_out           => s_data_out(10,45),
			out1               => s_out1(10,45),
			out2               => s_out2(10,45),
			lock_lower_row_out => s_locks_lower_out(10,45),
			lock_lower_row_in  => s_locks_lower_in(10,45),
			in1                => s_in1(10,45),
			in2                => s_in2(10,45),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(45)
		);
	s_in1(10,45)            <= s_out1(11,45);
	s_in2(10,45)            <= s_out2(11,46);
	s_locks_lower_in(10,45) <= s_locks_lower_out(11,45);

		normal_cell_10_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,46),
			fetch              => s_fetch(10,46),
			data_in            => s_data_in(10,46),
			data_out           => s_data_out(10,46),
			out1               => s_out1(10,46),
			out2               => s_out2(10,46),
			lock_lower_row_out => s_locks_lower_out(10,46),
			lock_lower_row_in  => s_locks_lower_in(10,46),
			in1                => s_in1(10,46),
			in2                => s_in2(10,46),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(46)
		);
	s_in1(10,46)            <= s_out1(11,46);
	s_in2(10,46)            <= s_out2(11,47);
	s_locks_lower_in(10,46) <= s_locks_lower_out(11,46);

		normal_cell_10_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,47),
			fetch              => s_fetch(10,47),
			data_in            => s_data_in(10,47),
			data_out           => s_data_out(10,47),
			out1               => s_out1(10,47),
			out2               => s_out2(10,47),
			lock_lower_row_out => s_locks_lower_out(10,47),
			lock_lower_row_in  => s_locks_lower_in(10,47),
			in1                => s_in1(10,47),
			in2                => s_in2(10,47),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(47)
		);
	s_in1(10,47)            <= s_out1(11,47);
	s_in2(10,47)            <= s_out2(11,48);
	s_locks_lower_in(10,47) <= s_locks_lower_out(11,47);

		normal_cell_10_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,48),
			fetch              => s_fetch(10,48),
			data_in            => s_data_in(10,48),
			data_out           => s_data_out(10,48),
			out1               => s_out1(10,48),
			out2               => s_out2(10,48),
			lock_lower_row_out => s_locks_lower_out(10,48),
			lock_lower_row_in  => s_locks_lower_in(10,48),
			in1                => s_in1(10,48),
			in2                => s_in2(10,48),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(48)
		);
	s_in1(10,48)            <= s_out1(11,48);
	s_in2(10,48)            <= s_out2(11,49);
	s_locks_lower_in(10,48) <= s_locks_lower_out(11,48);

		normal_cell_10_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,49),
			fetch              => s_fetch(10,49),
			data_in            => s_data_in(10,49),
			data_out           => s_data_out(10,49),
			out1               => s_out1(10,49),
			out2               => s_out2(10,49),
			lock_lower_row_out => s_locks_lower_out(10,49),
			lock_lower_row_in  => s_locks_lower_in(10,49),
			in1                => s_in1(10,49),
			in2                => s_in2(10,49),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(49)
		);
	s_in1(10,49)            <= s_out1(11,49);
	s_in2(10,49)            <= s_out2(11,50);
	s_locks_lower_in(10,49) <= s_locks_lower_out(11,49);

		normal_cell_10_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,50),
			fetch              => s_fetch(10,50),
			data_in            => s_data_in(10,50),
			data_out           => s_data_out(10,50),
			out1               => s_out1(10,50),
			out2               => s_out2(10,50),
			lock_lower_row_out => s_locks_lower_out(10,50),
			lock_lower_row_in  => s_locks_lower_in(10,50),
			in1                => s_in1(10,50),
			in2                => s_in2(10,50),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(50)
		);
	s_in1(10,50)            <= s_out1(11,50);
	s_in2(10,50)            <= s_out2(11,51);
	s_locks_lower_in(10,50) <= s_locks_lower_out(11,50);

		normal_cell_10_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,51),
			fetch              => s_fetch(10,51),
			data_in            => s_data_in(10,51),
			data_out           => s_data_out(10,51),
			out1               => s_out1(10,51),
			out2               => s_out2(10,51),
			lock_lower_row_out => s_locks_lower_out(10,51),
			lock_lower_row_in  => s_locks_lower_in(10,51),
			in1                => s_in1(10,51),
			in2                => s_in2(10,51),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(51)
		);
	s_in1(10,51)            <= s_out1(11,51);
	s_in2(10,51)            <= s_out2(11,52);
	s_locks_lower_in(10,51) <= s_locks_lower_out(11,51);

		normal_cell_10_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,52),
			fetch              => s_fetch(10,52),
			data_in            => s_data_in(10,52),
			data_out           => s_data_out(10,52),
			out1               => s_out1(10,52),
			out2               => s_out2(10,52),
			lock_lower_row_out => s_locks_lower_out(10,52),
			lock_lower_row_in  => s_locks_lower_in(10,52),
			in1                => s_in1(10,52),
			in2                => s_in2(10,52),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(52)
		);
	s_in1(10,52)            <= s_out1(11,52);
	s_in2(10,52)            <= s_out2(11,53);
	s_locks_lower_in(10,52) <= s_locks_lower_out(11,52);

		normal_cell_10_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,53),
			fetch              => s_fetch(10,53),
			data_in            => s_data_in(10,53),
			data_out           => s_data_out(10,53),
			out1               => s_out1(10,53),
			out2               => s_out2(10,53),
			lock_lower_row_out => s_locks_lower_out(10,53),
			lock_lower_row_in  => s_locks_lower_in(10,53),
			in1                => s_in1(10,53),
			in2                => s_in2(10,53),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(53)
		);
	s_in1(10,53)            <= s_out1(11,53);
	s_in2(10,53)            <= s_out2(11,54);
	s_locks_lower_in(10,53) <= s_locks_lower_out(11,53);

		normal_cell_10_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,54),
			fetch              => s_fetch(10,54),
			data_in            => s_data_in(10,54),
			data_out           => s_data_out(10,54),
			out1               => s_out1(10,54),
			out2               => s_out2(10,54),
			lock_lower_row_out => s_locks_lower_out(10,54),
			lock_lower_row_in  => s_locks_lower_in(10,54),
			in1                => s_in1(10,54),
			in2                => s_in2(10,54),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(54)
		);
	s_in1(10,54)            <= s_out1(11,54);
	s_in2(10,54)            <= s_out2(11,55);
	s_locks_lower_in(10,54) <= s_locks_lower_out(11,54);

		normal_cell_10_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,55),
			fetch              => s_fetch(10,55),
			data_in            => s_data_in(10,55),
			data_out           => s_data_out(10,55),
			out1               => s_out1(10,55),
			out2               => s_out2(10,55),
			lock_lower_row_out => s_locks_lower_out(10,55),
			lock_lower_row_in  => s_locks_lower_in(10,55),
			in1                => s_in1(10,55),
			in2                => s_in2(10,55),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(55)
		);
	s_in1(10,55)            <= s_out1(11,55);
	s_in2(10,55)            <= s_out2(11,56);
	s_locks_lower_in(10,55) <= s_locks_lower_out(11,55);

		normal_cell_10_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,56),
			fetch              => s_fetch(10,56),
			data_in            => s_data_in(10,56),
			data_out           => s_data_out(10,56),
			out1               => s_out1(10,56),
			out2               => s_out2(10,56),
			lock_lower_row_out => s_locks_lower_out(10,56),
			lock_lower_row_in  => s_locks_lower_in(10,56),
			in1                => s_in1(10,56),
			in2                => s_in2(10,56),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(56)
		);
	s_in1(10,56)            <= s_out1(11,56);
	s_in2(10,56)            <= s_out2(11,57);
	s_locks_lower_in(10,56) <= s_locks_lower_out(11,56);

		normal_cell_10_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,57),
			fetch              => s_fetch(10,57),
			data_in            => s_data_in(10,57),
			data_out           => s_data_out(10,57),
			out1               => s_out1(10,57),
			out2               => s_out2(10,57),
			lock_lower_row_out => s_locks_lower_out(10,57),
			lock_lower_row_in  => s_locks_lower_in(10,57),
			in1                => s_in1(10,57),
			in2                => s_in2(10,57),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(57)
		);
	s_in1(10,57)            <= s_out1(11,57);
	s_in2(10,57)            <= s_out2(11,58);
	s_locks_lower_in(10,57) <= s_locks_lower_out(11,57);

		normal_cell_10_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,58),
			fetch              => s_fetch(10,58),
			data_in            => s_data_in(10,58),
			data_out           => s_data_out(10,58),
			out1               => s_out1(10,58),
			out2               => s_out2(10,58),
			lock_lower_row_out => s_locks_lower_out(10,58),
			lock_lower_row_in  => s_locks_lower_in(10,58),
			in1                => s_in1(10,58),
			in2                => s_in2(10,58),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(58)
		);
	s_in1(10,58)            <= s_out1(11,58);
	s_in2(10,58)            <= s_out2(11,59);
	s_locks_lower_in(10,58) <= s_locks_lower_out(11,58);

		normal_cell_10_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,59),
			fetch              => s_fetch(10,59),
			data_in            => s_data_in(10,59),
			data_out           => s_data_out(10,59),
			out1               => s_out1(10,59),
			out2               => s_out2(10,59),
			lock_lower_row_out => s_locks_lower_out(10,59),
			lock_lower_row_in  => s_locks_lower_in(10,59),
			in1                => s_in1(10,59),
			in2                => s_in2(10,59),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(59)
		);
	s_in1(10,59)            <= s_out1(11,59);
	s_in2(10,59)            <= s_out2(11,60);
	s_locks_lower_in(10,59) <= s_locks_lower_out(11,59);

		last_col_cell_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(10,60),
			fetch              => s_fetch(10,60),
			data_in            => s_data_in(10,60),
			data_out           => s_data_out(10,60),
			out1               => s_out1(10,60),
			out2               => s_out2(10,60),
			lock_lower_row_out => s_locks_lower_out(10,60),
			lock_lower_row_in  => s_locks_lower_in(10,60),
			in1                => s_in1(10,60),
			in2                => (others => '0'),
			lock_row           => s_locks(10),
			piv_found          => s_piv_found,
			row_data           => s_row_data(10),
			col_data           => s_col_data(60)
		);
	s_in1(10,60)            <= s_out1(11,60);
	s_locks_lower_in(10,60) <= s_locks_lower_out(11,60);

		normal_cell_11_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,1),
			fetch              => s_fetch(11,1),
			data_in            => s_data_in(11,1),
			data_out           => s_data_out(11,1),
			out1               => s_out1(11,1),
			out2               => s_out2(11,1),
			lock_lower_row_out => s_locks_lower_out(11,1),
			lock_lower_row_in  => s_locks_lower_in(11,1),
			in1                => s_in1(11,1),
			in2                => s_in2(11,1),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(1)
		);
	s_in1(11,1)            <= s_out1(12,1);
	s_in2(11,1)            <= s_out2(12,2);
	s_locks_lower_in(11,1) <= s_locks_lower_out(12,1);

		normal_cell_11_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,2),
			fetch              => s_fetch(11,2),
			data_in            => s_data_in(11,2),
			data_out           => s_data_out(11,2),
			out1               => s_out1(11,2),
			out2               => s_out2(11,2),
			lock_lower_row_out => s_locks_lower_out(11,2),
			lock_lower_row_in  => s_locks_lower_in(11,2),
			in1                => s_in1(11,2),
			in2                => s_in2(11,2),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(2)
		);
	s_in1(11,2)            <= s_out1(12,2);
	s_in2(11,2)            <= s_out2(12,3);
	s_locks_lower_in(11,2) <= s_locks_lower_out(12,2);

		normal_cell_11_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,3),
			fetch              => s_fetch(11,3),
			data_in            => s_data_in(11,3),
			data_out           => s_data_out(11,3),
			out1               => s_out1(11,3),
			out2               => s_out2(11,3),
			lock_lower_row_out => s_locks_lower_out(11,3),
			lock_lower_row_in  => s_locks_lower_in(11,3),
			in1                => s_in1(11,3),
			in2                => s_in2(11,3),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(3)
		);
	s_in1(11,3)            <= s_out1(12,3);
	s_in2(11,3)            <= s_out2(12,4);
	s_locks_lower_in(11,3) <= s_locks_lower_out(12,3);

		normal_cell_11_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,4),
			fetch              => s_fetch(11,4),
			data_in            => s_data_in(11,4),
			data_out           => s_data_out(11,4),
			out1               => s_out1(11,4),
			out2               => s_out2(11,4),
			lock_lower_row_out => s_locks_lower_out(11,4),
			lock_lower_row_in  => s_locks_lower_in(11,4),
			in1                => s_in1(11,4),
			in2                => s_in2(11,4),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(4)
		);
	s_in1(11,4)            <= s_out1(12,4);
	s_in2(11,4)            <= s_out2(12,5);
	s_locks_lower_in(11,4) <= s_locks_lower_out(12,4);

		normal_cell_11_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,5),
			fetch              => s_fetch(11,5),
			data_in            => s_data_in(11,5),
			data_out           => s_data_out(11,5),
			out1               => s_out1(11,5),
			out2               => s_out2(11,5),
			lock_lower_row_out => s_locks_lower_out(11,5),
			lock_lower_row_in  => s_locks_lower_in(11,5),
			in1                => s_in1(11,5),
			in2                => s_in2(11,5),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(5)
		);
	s_in1(11,5)            <= s_out1(12,5);
	s_in2(11,5)            <= s_out2(12,6);
	s_locks_lower_in(11,5) <= s_locks_lower_out(12,5);

		normal_cell_11_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,6),
			fetch              => s_fetch(11,6),
			data_in            => s_data_in(11,6),
			data_out           => s_data_out(11,6),
			out1               => s_out1(11,6),
			out2               => s_out2(11,6),
			lock_lower_row_out => s_locks_lower_out(11,6),
			lock_lower_row_in  => s_locks_lower_in(11,6),
			in1                => s_in1(11,6),
			in2                => s_in2(11,6),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(6)
		);
	s_in1(11,6)            <= s_out1(12,6);
	s_in2(11,6)            <= s_out2(12,7);
	s_locks_lower_in(11,6) <= s_locks_lower_out(12,6);

		normal_cell_11_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,7),
			fetch              => s_fetch(11,7),
			data_in            => s_data_in(11,7),
			data_out           => s_data_out(11,7),
			out1               => s_out1(11,7),
			out2               => s_out2(11,7),
			lock_lower_row_out => s_locks_lower_out(11,7),
			lock_lower_row_in  => s_locks_lower_in(11,7),
			in1                => s_in1(11,7),
			in2                => s_in2(11,7),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(7)
		);
	s_in1(11,7)            <= s_out1(12,7);
	s_in2(11,7)            <= s_out2(12,8);
	s_locks_lower_in(11,7) <= s_locks_lower_out(12,7);

		normal_cell_11_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,8),
			fetch              => s_fetch(11,8),
			data_in            => s_data_in(11,8),
			data_out           => s_data_out(11,8),
			out1               => s_out1(11,8),
			out2               => s_out2(11,8),
			lock_lower_row_out => s_locks_lower_out(11,8),
			lock_lower_row_in  => s_locks_lower_in(11,8),
			in1                => s_in1(11,8),
			in2                => s_in2(11,8),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(8)
		);
	s_in1(11,8)            <= s_out1(12,8);
	s_in2(11,8)            <= s_out2(12,9);
	s_locks_lower_in(11,8) <= s_locks_lower_out(12,8);

		normal_cell_11_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,9),
			fetch              => s_fetch(11,9),
			data_in            => s_data_in(11,9),
			data_out           => s_data_out(11,9),
			out1               => s_out1(11,9),
			out2               => s_out2(11,9),
			lock_lower_row_out => s_locks_lower_out(11,9),
			lock_lower_row_in  => s_locks_lower_in(11,9),
			in1                => s_in1(11,9),
			in2                => s_in2(11,9),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(9)
		);
	s_in1(11,9)            <= s_out1(12,9);
	s_in2(11,9)            <= s_out2(12,10);
	s_locks_lower_in(11,9) <= s_locks_lower_out(12,9);

		normal_cell_11_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,10),
			fetch              => s_fetch(11,10),
			data_in            => s_data_in(11,10),
			data_out           => s_data_out(11,10),
			out1               => s_out1(11,10),
			out2               => s_out2(11,10),
			lock_lower_row_out => s_locks_lower_out(11,10),
			lock_lower_row_in  => s_locks_lower_in(11,10),
			in1                => s_in1(11,10),
			in2                => s_in2(11,10),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(10)
		);
	s_in1(11,10)            <= s_out1(12,10);
	s_in2(11,10)            <= s_out2(12,11);
	s_locks_lower_in(11,10) <= s_locks_lower_out(12,10);

		normal_cell_11_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,11),
			fetch              => s_fetch(11,11),
			data_in            => s_data_in(11,11),
			data_out           => s_data_out(11,11),
			out1               => s_out1(11,11),
			out2               => s_out2(11,11),
			lock_lower_row_out => s_locks_lower_out(11,11),
			lock_lower_row_in  => s_locks_lower_in(11,11),
			in1                => s_in1(11,11),
			in2                => s_in2(11,11),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(11)
		);
	s_in1(11,11)            <= s_out1(12,11);
	s_in2(11,11)            <= s_out2(12,12);
	s_locks_lower_in(11,11) <= s_locks_lower_out(12,11);

		normal_cell_11_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,12),
			fetch              => s_fetch(11,12),
			data_in            => s_data_in(11,12),
			data_out           => s_data_out(11,12),
			out1               => s_out1(11,12),
			out2               => s_out2(11,12),
			lock_lower_row_out => s_locks_lower_out(11,12),
			lock_lower_row_in  => s_locks_lower_in(11,12),
			in1                => s_in1(11,12),
			in2                => s_in2(11,12),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(12)
		);
	s_in1(11,12)            <= s_out1(12,12);
	s_in2(11,12)            <= s_out2(12,13);
	s_locks_lower_in(11,12) <= s_locks_lower_out(12,12);

		normal_cell_11_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,13),
			fetch              => s_fetch(11,13),
			data_in            => s_data_in(11,13),
			data_out           => s_data_out(11,13),
			out1               => s_out1(11,13),
			out2               => s_out2(11,13),
			lock_lower_row_out => s_locks_lower_out(11,13),
			lock_lower_row_in  => s_locks_lower_in(11,13),
			in1                => s_in1(11,13),
			in2                => s_in2(11,13),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(13)
		);
	s_in1(11,13)            <= s_out1(12,13);
	s_in2(11,13)            <= s_out2(12,14);
	s_locks_lower_in(11,13) <= s_locks_lower_out(12,13);

		normal_cell_11_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,14),
			fetch              => s_fetch(11,14),
			data_in            => s_data_in(11,14),
			data_out           => s_data_out(11,14),
			out1               => s_out1(11,14),
			out2               => s_out2(11,14),
			lock_lower_row_out => s_locks_lower_out(11,14),
			lock_lower_row_in  => s_locks_lower_in(11,14),
			in1                => s_in1(11,14),
			in2                => s_in2(11,14),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(14)
		);
	s_in1(11,14)            <= s_out1(12,14);
	s_in2(11,14)            <= s_out2(12,15);
	s_locks_lower_in(11,14) <= s_locks_lower_out(12,14);

		normal_cell_11_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,15),
			fetch              => s_fetch(11,15),
			data_in            => s_data_in(11,15),
			data_out           => s_data_out(11,15),
			out1               => s_out1(11,15),
			out2               => s_out2(11,15),
			lock_lower_row_out => s_locks_lower_out(11,15),
			lock_lower_row_in  => s_locks_lower_in(11,15),
			in1                => s_in1(11,15),
			in2                => s_in2(11,15),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(15)
		);
	s_in1(11,15)            <= s_out1(12,15);
	s_in2(11,15)            <= s_out2(12,16);
	s_locks_lower_in(11,15) <= s_locks_lower_out(12,15);

		normal_cell_11_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,16),
			fetch              => s_fetch(11,16),
			data_in            => s_data_in(11,16),
			data_out           => s_data_out(11,16),
			out1               => s_out1(11,16),
			out2               => s_out2(11,16),
			lock_lower_row_out => s_locks_lower_out(11,16),
			lock_lower_row_in  => s_locks_lower_in(11,16),
			in1                => s_in1(11,16),
			in2                => s_in2(11,16),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(16)
		);
	s_in1(11,16)            <= s_out1(12,16);
	s_in2(11,16)            <= s_out2(12,17);
	s_locks_lower_in(11,16) <= s_locks_lower_out(12,16);

		normal_cell_11_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,17),
			fetch              => s_fetch(11,17),
			data_in            => s_data_in(11,17),
			data_out           => s_data_out(11,17),
			out1               => s_out1(11,17),
			out2               => s_out2(11,17),
			lock_lower_row_out => s_locks_lower_out(11,17),
			lock_lower_row_in  => s_locks_lower_in(11,17),
			in1                => s_in1(11,17),
			in2                => s_in2(11,17),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(17)
		);
	s_in1(11,17)            <= s_out1(12,17);
	s_in2(11,17)            <= s_out2(12,18);
	s_locks_lower_in(11,17) <= s_locks_lower_out(12,17);

		normal_cell_11_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,18),
			fetch              => s_fetch(11,18),
			data_in            => s_data_in(11,18),
			data_out           => s_data_out(11,18),
			out1               => s_out1(11,18),
			out2               => s_out2(11,18),
			lock_lower_row_out => s_locks_lower_out(11,18),
			lock_lower_row_in  => s_locks_lower_in(11,18),
			in1                => s_in1(11,18),
			in2                => s_in2(11,18),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(18)
		);
	s_in1(11,18)            <= s_out1(12,18);
	s_in2(11,18)            <= s_out2(12,19);
	s_locks_lower_in(11,18) <= s_locks_lower_out(12,18);

		normal_cell_11_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,19),
			fetch              => s_fetch(11,19),
			data_in            => s_data_in(11,19),
			data_out           => s_data_out(11,19),
			out1               => s_out1(11,19),
			out2               => s_out2(11,19),
			lock_lower_row_out => s_locks_lower_out(11,19),
			lock_lower_row_in  => s_locks_lower_in(11,19),
			in1                => s_in1(11,19),
			in2                => s_in2(11,19),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(19)
		);
	s_in1(11,19)            <= s_out1(12,19);
	s_in2(11,19)            <= s_out2(12,20);
	s_locks_lower_in(11,19) <= s_locks_lower_out(12,19);

		normal_cell_11_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,20),
			fetch              => s_fetch(11,20),
			data_in            => s_data_in(11,20),
			data_out           => s_data_out(11,20),
			out1               => s_out1(11,20),
			out2               => s_out2(11,20),
			lock_lower_row_out => s_locks_lower_out(11,20),
			lock_lower_row_in  => s_locks_lower_in(11,20),
			in1                => s_in1(11,20),
			in2                => s_in2(11,20),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(20)
		);
	s_in1(11,20)            <= s_out1(12,20);
	s_in2(11,20)            <= s_out2(12,21);
	s_locks_lower_in(11,20) <= s_locks_lower_out(12,20);

		normal_cell_11_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,21),
			fetch              => s_fetch(11,21),
			data_in            => s_data_in(11,21),
			data_out           => s_data_out(11,21),
			out1               => s_out1(11,21),
			out2               => s_out2(11,21),
			lock_lower_row_out => s_locks_lower_out(11,21),
			lock_lower_row_in  => s_locks_lower_in(11,21),
			in1                => s_in1(11,21),
			in2                => s_in2(11,21),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(21)
		);
	s_in1(11,21)            <= s_out1(12,21);
	s_in2(11,21)            <= s_out2(12,22);
	s_locks_lower_in(11,21) <= s_locks_lower_out(12,21);

		normal_cell_11_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,22),
			fetch              => s_fetch(11,22),
			data_in            => s_data_in(11,22),
			data_out           => s_data_out(11,22),
			out1               => s_out1(11,22),
			out2               => s_out2(11,22),
			lock_lower_row_out => s_locks_lower_out(11,22),
			lock_lower_row_in  => s_locks_lower_in(11,22),
			in1                => s_in1(11,22),
			in2                => s_in2(11,22),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(22)
		);
	s_in1(11,22)            <= s_out1(12,22);
	s_in2(11,22)            <= s_out2(12,23);
	s_locks_lower_in(11,22) <= s_locks_lower_out(12,22);

		normal_cell_11_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,23),
			fetch              => s_fetch(11,23),
			data_in            => s_data_in(11,23),
			data_out           => s_data_out(11,23),
			out1               => s_out1(11,23),
			out2               => s_out2(11,23),
			lock_lower_row_out => s_locks_lower_out(11,23),
			lock_lower_row_in  => s_locks_lower_in(11,23),
			in1                => s_in1(11,23),
			in2                => s_in2(11,23),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(23)
		);
	s_in1(11,23)            <= s_out1(12,23);
	s_in2(11,23)            <= s_out2(12,24);
	s_locks_lower_in(11,23) <= s_locks_lower_out(12,23);

		normal_cell_11_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,24),
			fetch              => s_fetch(11,24),
			data_in            => s_data_in(11,24),
			data_out           => s_data_out(11,24),
			out1               => s_out1(11,24),
			out2               => s_out2(11,24),
			lock_lower_row_out => s_locks_lower_out(11,24),
			lock_lower_row_in  => s_locks_lower_in(11,24),
			in1                => s_in1(11,24),
			in2                => s_in2(11,24),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(24)
		);
	s_in1(11,24)            <= s_out1(12,24);
	s_in2(11,24)            <= s_out2(12,25);
	s_locks_lower_in(11,24) <= s_locks_lower_out(12,24);

		normal_cell_11_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,25),
			fetch              => s_fetch(11,25),
			data_in            => s_data_in(11,25),
			data_out           => s_data_out(11,25),
			out1               => s_out1(11,25),
			out2               => s_out2(11,25),
			lock_lower_row_out => s_locks_lower_out(11,25),
			lock_lower_row_in  => s_locks_lower_in(11,25),
			in1                => s_in1(11,25),
			in2                => s_in2(11,25),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(25)
		);
	s_in1(11,25)            <= s_out1(12,25);
	s_in2(11,25)            <= s_out2(12,26);
	s_locks_lower_in(11,25) <= s_locks_lower_out(12,25);

		normal_cell_11_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,26),
			fetch              => s_fetch(11,26),
			data_in            => s_data_in(11,26),
			data_out           => s_data_out(11,26),
			out1               => s_out1(11,26),
			out2               => s_out2(11,26),
			lock_lower_row_out => s_locks_lower_out(11,26),
			lock_lower_row_in  => s_locks_lower_in(11,26),
			in1                => s_in1(11,26),
			in2                => s_in2(11,26),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(26)
		);
	s_in1(11,26)            <= s_out1(12,26);
	s_in2(11,26)            <= s_out2(12,27);
	s_locks_lower_in(11,26) <= s_locks_lower_out(12,26);

		normal_cell_11_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,27),
			fetch              => s_fetch(11,27),
			data_in            => s_data_in(11,27),
			data_out           => s_data_out(11,27),
			out1               => s_out1(11,27),
			out2               => s_out2(11,27),
			lock_lower_row_out => s_locks_lower_out(11,27),
			lock_lower_row_in  => s_locks_lower_in(11,27),
			in1                => s_in1(11,27),
			in2                => s_in2(11,27),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(27)
		);
	s_in1(11,27)            <= s_out1(12,27);
	s_in2(11,27)            <= s_out2(12,28);
	s_locks_lower_in(11,27) <= s_locks_lower_out(12,27);

		normal_cell_11_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,28),
			fetch              => s_fetch(11,28),
			data_in            => s_data_in(11,28),
			data_out           => s_data_out(11,28),
			out1               => s_out1(11,28),
			out2               => s_out2(11,28),
			lock_lower_row_out => s_locks_lower_out(11,28),
			lock_lower_row_in  => s_locks_lower_in(11,28),
			in1                => s_in1(11,28),
			in2                => s_in2(11,28),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(28)
		);
	s_in1(11,28)            <= s_out1(12,28);
	s_in2(11,28)            <= s_out2(12,29);
	s_locks_lower_in(11,28) <= s_locks_lower_out(12,28);

		normal_cell_11_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,29),
			fetch              => s_fetch(11,29),
			data_in            => s_data_in(11,29),
			data_out           => s_data_out(11,29),
			out1               => s_out1(11,29),
			out2               => s_out2(11,29),
			lock_lower_row_out => s_locks_lower_out(11,29),
			lock_lower_row_in  => s_locks_lower_in(11,29),
			in1                => s_in1(11,29),
			in2                => s_in2(11,29),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(29)
		);
	s_in1(11,29)            <= s_out1(12,29);
	s_in2(11,29)            <= s_out2(12,30);
	s_locks_lower_in(11,29) <= s_locks_lower_out(12,29);

		normal_cell_11_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,30),
			fetch              => s_fetch(11,30),
			data_in            => s_data_in(11,30),
			data_out           => s_data_out(11,30),
			out1               => s_out1(11,30),
			out2               => s_out2(11,30),
			lock_lower_row_out => s_locks_lower_out(11,30),
			lock_lower_row_in  => s_locks_lower_in(11,30),
			in1                => s_in1(11,30),
			in2                => s_in2(11,30),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(30)
		);
	s_in1(11,30)            <= s_out1(12,30);
	s_in2(11,30)            <= s_out2(12,31);
	s_locks_lower_in(11,30) <= s_locks_lower_out(12,30);

		normal_cell_11_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,31),
			fetch              => s_fetch(11,31),
			data_in            => s_data_in(11,31),
			data_out           => s_data_out(11,31),
			out1               => s_out1(11,31),
			out2               => s_out2(11,31),
			lock_lower_row_out => s_locks_lower_out(11,31),
			lock_lower_row_in  => s_locks_lower_in(11,31),
			in1                => s_in1(11,31),
			in2                => s_in2(11,31),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(31)
		);
	s_in1(11,31)            <= s_out1(12,31);
	s_in2(11,31)            <= s_out2(12,32);
	s_locks_lower_in(11,31) <= s_locks_lower_out(12,31);

		normal_cell_11_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,32),
			fetch              => s_fetch(11,32),
			data_in            => s_data_in(11,32),
			data_out           => s_data_out(11,32),
			out1               => s_out1(11,32),
			out2               => s_out2(11,32),
			lock_lower_row_out => s_locks_lower_out(11,32),
			lock_lower_row_in  => s_locks_lower_in(11,32),
			in1                => s_in1(11,32),
			in2                => s_in2(11,32),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(32)
		);
	s_in1(11,32)            <= s_out1(12,32);
	s_in2(11,32)            <= s_out2(12,33);
	s_locks_lower_in(11,32) <= s_locks_lower_out(12,32);

		normal_cell_11_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,33),
			fetch              => s_fetch(11,33),
			data_in            => s_data_in(11,33),
			data_out           => s_data_out(11,33),
			out1               => s_out1(11,33),
			out2               => s_out2(11,33),
			lock_lower_row_out => s_locks_lower_out(11,33),
			lock_lower_row_in  => s_locks_lower_in(11,33),
			in1                => s_in1(11,33),
			in2                => s_in2(11,33),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(33)
		);
	s_in1(11,33)            <= s_out1(12,33);
	s_in2(11,33)            <= s_out2(12,34);
	s_locks_lower_in(11,33) <= s_locks_lower_out(12,33);

		normal_cell_11_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,34),
			fetch              => s_fetch(11,34),
			data_in            => s_data_in(11,34),
			data_out           => s_data_out(11,34),
			out1               => s_out1(11,34),
			out2               => s_out2(11,34),
			lock_lower_row_out => s_locks_lower_out(11,34),
			lock_lower_row_in  => s_locks_lower_in(11,34),
			in1                => s_in1(11,34),
			in2                => s_in2(11,34),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(34)
		);
	s_in1(11,34)            <= s_out1(12,34);
	s_in2(11,34)            <= s_out2(12,35);
	s_locks_lower_in(11,34) <= s_locks_lower_out(12,34);

		normal_cell_11_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,35),
			fetch              => s_fetch(11,35),
			data_in            => s_data_in(11,35),
			data_out           => s_data_out(11,35),
			out1               => s_out1(11,35),
			out2               => s_out2(11,35),
			lock_lower_row_out => s_locks_lower_out(11,35),
			lock_lower_row_in  => s_locks_lower_in(11,35),
			in1                => s_in1(11,35),
			in2                => s_in2(11,35),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(35)
		);
	s_in1(11,35)            <= s_out1(12,35);
	s_in2(11,35)            <= s_out2(12,36);
	s_locks_lower_in(11,35) <= s_locks_lower_out(12,35);

		normal_cell_11_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,36),
			fetch              => s_fetch(11,36),
			data_in            => s_data_in(11,36),
			data_out           => s_data_out(11,36),
			out1               => s_out1(11,36),
			out2               => s_out2(11,36),
			lock_lower_row_out => s_locks_lower_out(11,36),
			lock_lower_row_in  => s_locks_lower_in(11,36),
			in1                => s_in1(11,36),
			in2                => s_in2(11,36),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(36)
		);
	s_in1(11,36)            <= s_out1(12,36);
	s_in2(11,36)            <= s_out2(12,37);
	s_locks_lower_in(11,36) <= s_locks_lower_out(12,36);

		normal_cell_11_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,37),
			fetch              => s_fetch(11,37),
			data_in            => s_data_in(11,37),
			data_out           => s_data_out(11,37),
			out1               => s_out1(11,37),
			out2               => s_out2(11,37),
			lock_lower_row_out => s_locks_lower_out(11,37),
			lock_lower_row_in  => s_locks_lower_in(11,37),
			in1                => s_in1(11,37),
			in2                => s_in2(11,37),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(37)
		);
	s_in1(11,37)            <= s_out1(12,37);
	s_in2(11,37)            <= s_out2(12,38);
	s_locks_lower_in(11,37) <= s_locks_lower_out(12,37);

		normal_cell_11_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,38),
			fetch              => s_fetch(11,38),
			data_in            => s_data_in(11,38),
			data_out           => s_data_out(11,38),
			out1               => s_out1(11,38),
			out2               => s_out2(11,38),
			lock_lower_row_out => s_locks_lower_out(11,38),
			lock_lower_row_in  => s_locks_lower_in(11,38),
			in1                => s_in1(11,38),
			in2                => s_in2(11,38),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(38)
		);
	s_in1(11,38)            <= s_out1(12,38);
	s_in2(11,38)            <= s_out2(12,39);
	s_locks_lower_in(11,38) <= s_locks_lower_out(12,38);

		normal_cell_11_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,39),
			fetch              => s_fetch(11,39),
			data_in            => s_data_in(11,39),
			data_out           => s_data_out(11,39),
			out1               => s_out1(11,39),
			out2               => s_out2(11,39),
			lock_lower_row_out => s_locks_lower_out(11,39),
			lock_lower_row_in  => s_locks_lower_in(11,39),
			in1                => s_in1(11,39),
			in2                => s_in2(11,39),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(39)
		);
	s_in1(11,39)            <= s_out1(12,39);
	s_in2(11,39)            <= s_out2(12,40);
	s_locks_lower_in(11,39) <= s_locks_lower_out(12,39);

		normal_cell_11_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,40),
			fetch              => s_fetch(11,40),
			data_in            => s_data_in(11,40),
			data_out           => s_data_out(11,40),
			out1               => s_out1(11,40),
			out2               => s_out2(11,40),
			lock_lower_row_out => s_locks_lower_out(11,40),
			lock_lower_row_in  => s_locks_lower_in(11,40),
			in1                => s_in1(11,40),
			in2                => s_in2(11,40),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(40)
		);
	s_in1(11,40)            <= s_out1(12,40);
	s_in2(11,40)            <= s_out2(12,41);
	s_locks_lower_in(11,40) <= s_locks_lower_out(12,40);

		normal_cell_11_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,41),
			fetch              => s_fetch(11,41),
			data_in            => s_data_in(11,41),
			data_out           => s_data_out(11,41),
			out1               => s_out1(11,41),
			out2               => s_out2(11,41),
			lock_lower_row_out => s_locks_lower_out(11,41),
			lock_lower_row_in  => s_locks_lower_in(11,41),
			in1                => s_in1(11,41),
			in2                => s_in2(11,41),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(41)
		);
	s_in1(11,41)            <= s_out1(12,41);
	s_in2(11,41)            <= s_out2(12,42);
	s_locks_lower_in(11,41) <= s_locks_lower_out(12,41);

		normal_cell_11_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,42),
			fetch              => s_fetch(11,42),
			data_in            => s_data_in(11,42),
			data_out           => s_data_out(11,42),
			out1               => s_out1(11,42),
			out2               => s_out2(11,42),
			lock_lower_row_out => s_locks_lower_out(11,42),
			lock_lower_row_in  => s_locks_lower_in(11,42),
			in1                => s_in1(11,42),
			in2                => s_in2(11,42),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(42)
		);
	s_in1(11,42)            <= s_out1(12,42);
	s_in2(11,42)            <= s_out2(12,43);
	s_locks_lower_in(11,42) <= s_locks_lower_out(12,42);

		normal_cell_11_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,43),
			fetch              => s_fetch(11,43),
			data_in            => s_data_in(11,43),
			data_out           => s_data_out(11,43),
			out1               => s_out1(11,43),
			out2               => s_out2(11,43),
			lock_lower_row_out => s_locks_lower_out(11,43),
			lock_lower_row_in  => s_locks_lower_in(11,43),
			in1                => s_in1(11,43),
			in2                => s_in2(11,43),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(43)
		);
	s_in1(11,43)            <= s_out1(12,43);
	s_in2(11,43)            <= s_out2(12,44);
	s_locks_lower_in(11,43) <= s_locks_lower_out(12,43);

		normal_cell_11_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,44),
			fetch              => s_fetch(11,44),
			data_in            => s_data_in(11,44),
			data_out           => s_data_out(11,44),
			out1               => s_out1(11,44),
			out2               => s_out2(11,44),
			lock_lower_row_out => s_locks_lower_out(11,44),
			lock_lower_row_in  => s_locks_lower_in(11,44),
			in1                => s_in1(11,44),
			in2                => s_in2(11,44),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(44)
		);
	s_in1(11,44)            <= s_out1(12,44);
	s_in2(11,44)            <= s_out2(12,45);
	s_locks_lower_in(11,44) <= s_locks_lower_out(12,44);

		normal_cell_11_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,45),
			fetch              => s_fetch(11,45),
			data_in            => s_data_in(11,45),
			data_out           => s_data_out(11,45),
			out1               => s_out1(11,45),
			out2               => s_out2(11,45),
			lock_lower_row_out => s_locks_lower_out(11,45),
			lock_lower_row_in  => s_locks_lower_in(11,45),
			in1                => s_in1(11,45),
			in2                => s_in2(11,45),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(45)
		);
	s_in1(11,45)            <= s_out1(12,45);
	s_in2(11,45)            <= s_out2(12,46);
	s_locks_lower_in(11,45) <= s_locks_lower_out(12,45);

		normal_cell_11_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,46),
			fetch              => s_fetch(11,46),
			data_in            => s_data_in(11,46),
			data_out           => s_data_out(11,46),
			out1               => s_out1(11,46),
			out2               => s_out2(11,46),
			lock_lower_row_out => s_locks_lower_out(11,46),
			lock_lower_row_in  => s_locks_lower_in(11,46),
			in1                => s_in1(11,46),
			in2                => s_in2(11,46),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(46)
		);
	s_in1(11,46)            <= s_out1(12,46);
	s_in2(11,46)            <= s_out2(12,47);
	s_locks_lower_in(11,46) <= s_locks_lower_out(12,46);

		normal_cell_11_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,47),
			fetch              => s_fetch(11,47),
			data_in            => s_data_in(11,47),
			data_out           => s_data_out(11,47),
			out1               => s_out1(11,47),
			out2               => s_out2(11,47),
			lock_lower_row_out => s_locks_lower_out(11,47),
			lock_lower_row_in  => s_locks_lower_in(11,47),
			in1                => s_in1(11,47),
			in2                => s_in2(11,47),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(47)
		);
	s_in1(11,47)            <= s_out1(12,47);
	s_in2(11,47)            <= s_out2(12,48);
	s_locks_lower_in(11,47) <= s_locks_lower_out(12,47);

		normal_cell_11_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,48),
			fetch              => s_fetch(11,48),
			data_in            => s_data_in(11,48),
			data_out           => s_data_out(11,48),
			out1               => s_out1(11,48),
			out2               => s_out2(11,48),
			lock_lower_row_out => s_locks_lower_out(11,48),
			lock_lower_row_in  => s_locks_lower_in(11,48),
			in1                => s_in1(11,48),
			in2                => s_in2(11,48),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(48)
		);
	s_in1(11,48)            <= s_out1(12,48);
	s_in2(11,48)            <= s_out2(12,49);
	s_locks_lower_in(11,48) <= s_locks_lower_out(12,48);

		normal_cell_11_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,49),
			fetch              => s_fetch(11,49),
			data_in            => s_data_in(11,49),
			data_out           => s_data_out(11,49),
			out1               => s_out1(11,49),
			out2               => s_out2(11,49),
			lock_lower_row_out => s_locks_lower_out(11,49),
			lock_lower_row_in  => s_locks_lower_in(11,49),
			in1                => s_in1(11,49),
			in2                => s_in2(11,49),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(49)
		);
	s_in1(11,49)            <= s_out1(12,49);
	s_in2(11,49)            <= s_out2(12,50);
	s_locks_lower_in(11,49) <= s_locks_lower_out(12,49);

		normal_cell_11_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,50),
			fetch              => s_fetch(11,50),
			data_in            => s_data_in(11,50),
			data_out           => s_data_out(11,50),
			out1               => s_out1(11,50),
			out2               => s_out2(11,50),
			lock_lower_row_out => s_locks_lower_out(11,50),
			lock_lower_row_in  => s_locks_lower_in(11,50),
			in1                => s_in1(11,50),
			in2                => s_in2(11,50),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(50)
		);
	s_in1(11,50)            <= s_out1(12,50);
	s_in2(11,50)            <= s_out2(12,51);
	s_locks_lower_in(11,50) <= s_locks_lower_out(12,50);

		normal_cell_11_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,51),
			fetch              => s_fetch(11,51),
			data_in            => s_data_in(11,51),
			data_out           => s_data_out(11,51),
			out1               => s_out1(11,51),
			out2               => s_out2(11,51),
			lock_lower_row_out => s_locks_lower_out(11,51),
			lock_lower_row_in  => s_locks_lower_in(11,51),
			in1                => s_in1(11,51),
			in2                => s_in2(11,51),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(51)
		);
	s_in1(11,51)            <= s_out1(12,51);
	s_in2(11,51)            <= s_out2(12,52);
	s_locks_lower_in(11,51) <= s_locks_lower_out(12,51);

		normal_cell_11_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,52),
			fetch              => s_fetch(11,52),
			data_in            => s_data_in(11,52),
			data_out           => s_data_out(11,52),
			out1               => s_out1(11,52),
			out2               => s_out2(11,52),
			lock_lower_row_out => s_locks_lower_out(11,52),
			lock_lower_row_in  => s_locks_lower_in(11,52),
			in1                => s_in1(11,52),
			in2                => s_in2(11,52),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(52)
		);
	s_in1(11,52)            <= s_out1(12,52);
	s_in2(11,52)            <= s_out2(12,53);
	s_locks_lower_in(11,52) <= s_locks_lower_out(12,52);

		normal_cell_11_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,53),
			fetch              => s_fetch(11,53),
			data_in            => s_data_in(11,53),
			data_out           => s_data_out(11,53),
			out1               => s_out1(11,53),
			out2               => s_out2(11,53),
			lock_lower_row_out => s_locks_lower_out(11,53),
			lock_lower_row_in  => s_locks_lower_in(11,53),
			in1                => s_in1(11,53),
			in2                => s_in2(11,53),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(53)
		);
	s_in1(11,53)            <= s_out1(12,53);
	s_in2(11,53)            <= s_out2(12,54);
	s_locks_lower_in(11,53) <= s_locks_lower_out(12,53);

		normal_cell_11_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,54),
			fetch              => s_fetch(11,54),
			data_in            => s_data_in(11,54),
			data_out           => s_data_out(11,54),
			out1               => s_out1(11,54),
			out2               => s_out2(11,54),
			lock_lower_row_out => s_locks_lower_out(11,54),
			lock_lower_row_in  => s_locks_lower_in(11,54),
			in1                => s_in1(11,54),
			in2                => s_in2(11,54),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(54)
		);
	s_in1(11,54)            <= s_out1(12,54);
	s_in2(11,54)            <= s_out2(12,55);
	s_locks_lower_in(11,54) <= s_locks_lower_out(12,54);

		normal_cell_11_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,55),
			fetch              => s_fetch(11,55),
			data_in            => s_data_in(11,55),
			data_out           => s_data_out(11,55),
			out1               => s_out1(11,55),
			out2               => s_out2(11,55),
			lock_lower_row_out => s_locks_lower_out(11,55),
			lock_lower_row_in  => s_locks_lower_in(11,55),
			in1                => s_in1(11,55),
			in2                => s_in2(11,55),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(55)
		);
	s_in1(11,55)            <= s_out1(12,55);
	s_in2(11,55)            <= s_out2(12,56);
	s_locks_lower_in(11,55) <= s_locks_lower_out(12,55);

		normal_cell_11_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,56),
			fetch              => s_fetch(11,56),
			data_in            => s_data_in(11,56),
			data_out           => s_data_out(11,56),
			out1               => s_out1(11,56),
			out2               => s_out2(11,56),
			lock_lower_row_out => s_locks_lower_out(11,56),
			lock_lower_row_in  => s_locks_lower_in(11,56),
			in1                => s_in1(11,56),
			in2                => s_in2(11,56),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(56)
		);
	s_in1(11,56)            <= s_out1(12,56);
	s_in2(11,56)            <= s_out2(12,57);
	s_locks_lower_in(11,56) <= s_locks_lower_out(12,56);

		normal_cell_11_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,57),
			fetch              => s_fetch(11,57),
			data_in            => s_data_in(11,57),
			data_out           => s_data_out(11,57),
			out1               => s_out1(11,57),
			out2               => s_out2(11,57),
			lock_lower_row_out => s_locks_lower_out(11,57),
			lock_lower_row_in  => s_locks_lower_in(11,57),
			in1                => s_in1(11,57),
			in2                => s_in2(11,57),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(57)
		);
	s_in1(11,57)            <= s_out1(12,57);
	s_in2(11,57)            <= s_out2(12,58);
	s_locks_lower_in(11,57) <= s_locks_lower_out(12,57);

		normal_cell_11_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,58),
			fetch              => s_fetch(11,58),
			data_in            => s_data_in(11,58),
			data_out           => s_data_out(11,58),
			out1               => s_out1(11,58),
			out2               => s_out2(11,58),
			lock_lower_row_out => s_locks_lower_out(11,58),
			lock_lower_row_in  => s_locks_lower_in(11,58),
			in1                => s_in1(11,58),
			in2                => s_in2(11,58),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(58)
		);
	s_in1(11,58)            <= s_out1(12,58);
	s_in2(11,58)            <= s_out2(12,59);
	s_locks_lower_in(11,58) <= s_locks_lower_out(12,58);

		normal_cell_11_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,59),
			fetch              => s_fetch(11,59),
			data_in            => s_data_in(11,59),
			data_out           => s_data_out(11,59),
			out1               => s_out1(11,59),
			out2               => s_out2(11,59),
			lock_lower_row_out => s_locks_lower_out(11,59),
			lock_lower_row_in  => s_locks_lower_in(11,59),
			in1                => s_in1(11,59),
			in2                => s_in2(11,59),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(59)
		);
	s_in1(11,59)            <= s_out1(12,59);
	s_in2(11,59)            <= s_out2(12,60);
	s_locks_lower_in(11,59) <= s_locks_lower_out(12,59);

		last_col_cell_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(11,60),
			fetch              => s_fetch(11,60),
			data_in            => s_data_in(11,60),
			data_out           => s_data_out(11,60),
			out1               => s_out1(11,60),
			out2               => s_out2(11,60),
			lock_lower_row_out => s_locks_lower_out(11,60),
			lock_lower_row_in  => s_locks_lower_in(11,60),
			in1                => s_in1(11,60),
			in2                => (others => '0'),
			lock_row           => s_locks(11),
			piv_found          => s_piv_found,
			row_data           => s_row_data(11),
			col_data           => s_col_data(60)
		);
	s_in1(11,60)            <= s_out1(12,60);
	s_locks_lower_in(11,60) <= s_locks_lower_out(12,60);

		normal_cell_12_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,1),
			fetch              => s_fetch(12,1),
			data_in            => s_data_in(12,1),
			data_out           => s_data_out(12,1),
			out1               => s_out1(12,1),
			out2               => s_out2(12,1),
			lock_lower_row_out => s_locks_lower_out(12,1),
			lock_lower_row_in  => s_locks_lower_in(12,1),
			in1                => s_in1(12,1),
			in2                => s_in2(12,1),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(1)
		);
	s_in1(12,1)            <= s_out1(13,1);
	s_in2(12,1)            <= s_out2(13,2);
	s_locks_lower_in(12,1) <= s_locks_lower_out(13,1);

		normal_cell_12_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,2),
			fetch              => s_fetch(12,2),
			data_in            => s_data_in(12,2),
			data_out           => s_data_out(12,2),
			out1               => s_out1(12,2),
			out2               => s_out2(12,2),
			lock_lower_row_out => s_locks_lower_out(12,2),
			lock_lower_row_in  => s_locks_lower_in(12,2),
			in1                => s_in1(12,2),
			in2                => s_in2(12,2),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(2)
		);
	s_in1(12,2)            <= s_out1(13,2);
	s_in2(12,2)            <= s_out2(13,3);
	s_locks_lower_in(12,2) <= s_locks_lower_out(13,2);

		normal_cell_12_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,3),
			fetch              => s_fetch(12,3),
			data_in            => s_data_in(12,3),
			data_out           => s_data_out(12,3),
			out1               => s_out1(12,3),
			out2               => s_out2(12,3),
			lock_lower_row_out => s_locks_lower_out(12,3),
			lock_lower_row_in  => s_locks_lower_in(12,3),
			in1                => s_in1(12,3),
			in2                => s_in2(12,3),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(3)
		);
	s_in1(12,3)            <= s_out1(13,3);
	s_in2(12,3)            <= s_out2(13,4);
	s_locks_lower_in(12,3) <= s_locks_lower_out(13,3);

		normal_cell_12_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,4),
			fetch              => s_fetch(12,4),
			data_in            => s_data_in(12,4),
			data_out           => s_data_out(12,4),
			out1               => s_out1(12,4),
			out2               => s_out2(12,4),
			lock_lower_row_out => s_locks_lower_out(12,4),
			lock_lower_row_in  => s_locks_lower_in(12,4),
			in1                => s_in1(12,4),
			in2                => s_in2(12,4),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(4)
		);
	s_in1(12,4)            <= s_out1(13,4);
	s_in2(12,4)            <= s_out2(13,5);
	s_locks_lower_in(12,4) <= s_locks_lower_out(13,4);

		normal_cell_12_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,5),
			fetch              => s_fetch(12,5),
			data_in            => s_data_in(12,5),
			data_out           => s_data_out(12,5),
			out1               => s_out1(12,5),
			out2               => s_out2(12,5),
			lock_lower_row_out => s_locks_lower_out(12,5),
			lock_lower_row_in  => s_locks_lower_in(12,5),
			in1                => s_in1(12,5),
			in2                => s_in2(12,5),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(5)
		);
	s_in1(12,5)            <= s_out1(13,5);
	s_in2(12,5)            <= s_out2(13,6);
	s_locks_lower_in(12,5) <= s_locks_lower_out(13,5);

		normal_cell_12_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,6),
			fetch              => s_fetch(12,6),
			data_in            => s_data_in(12,6),
			data_out           => s_data_out(12,6),
			out1               => s_out1(12,6),
			out2               => s_out2(12,6),
			lock_lower_row_out => s_locks_lower_out(12,6),
			lock_lower_row_in  => s_locks_lower_in(12,6),
			in1                => s_in1(12,6),
			in2                => s_in2(12,6),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(6)
		);
	s_in1(12,6)            <= s_out1(13,6);
	s_in2(12,6)            <= s_out2(13,7);
	s_locks_lower_in(12,6) <= s_locks_lower_out(13,6);

		normal_cell_12_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,7),
			fetch              => s_fetch(12,7),
			data_in            => s_data_in(12,7),
			data_out           => s_data_out(12,7),
			out1               => s_out1(12,7),
			out2               => s_out2(12,7),
			lock_lower_row_out => s_locks_lower_out(12,7),
			lock_lower_row_in  => s_locks_lower_in(12,7),
			in1                => s_in1(12,7),
			in2                => s_in2(12,7),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(7)
		);
	s_in1(12,7)            <= s_out1(13,7);
	s_in2(12,7)            <= s_out2(13,8);
	s_locks_lower_in(12,7) <= s_locks_lower_out(13,7);

		normal_cell_12_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,8),
			fetch              => s_fetch(12,8),
			data_in            => s_data_in(12,8),
			data_out           => s_data_out(12,8),
			out1               => s_out1(12,8),
			out2               => s_out2(12,8),
			lock_lower_row_out => s_locks_lower_out(12,8),
			lock_lower_row_in  => s_locks_lower_in(12,8),
			in1                => s_in1(12,8),
			in2                => s_in2(12,8),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(8)
		);
	s_in1(12,8)            <= s_out1(13,8);
	s_in2(12,8)            <= s_out2(13,9);
	s_locks_lower_in(12,8) <= s_locks_lower_out(13,8);

		normal_cell_12_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,9),
			fetch              => s_fetch(12,9),
			data_in            => s_data_in(12,9),
			data_out           => s_data_out(12,9),
			out1               => s_out1(12,9),
			out2               => s_out2(12,9),
			lock_lower_row_out => s_locks_lower_out(12,9),
			lock_lower_row_in  => s_locks_lower_in(12,9),
			in1                => s_in1(12,9),
			in2                => s_in2(12,9),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(9)
		);
	s_in1(12,9)            <= s_out1(13,9);
	s_in2(12,9)            <= s_out2(13,10);
	s_locks_lower_in(12,9) <= s_locks_lower_out(13,9);

		normal_cell_12_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,10),
			fetch              => s_fetch(12,10),
			data_in            => s_data_in(12,10),
			data_out           => s_data_out(12,10),
			out1               => s_out1(12,10),
			out2               => s_out2(12,10),
			lock_lower_row_out => s_locks_lower_out(12,10),
			lock_lower_row_in  => s_locks_lower_in(12,10),
			in1                => s_in1(12,10),
			in2                => s_in2(12,10),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(10)
		);
	s_in1(12,10)            <= s_out1(13,10);
	s_in2(12,10)            <= s_out2(13,11);
	s_locks_lower_in(12,10) <= s_locks_lower_out(13,10);

		normal_cell_12_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,11),
			fetch              => s_fetch(12,11),
			data_in            => s_data_in(12,11),
			data_out           => s_data_out(12,11),
			out1               => s_out1(12,11),
			out2               => s_out2(12,11),
			lock_lower_row_out => s_locks_lower_out(12,11),
			lock_lower_row_in  => s_locks_lower_in(12,11),
			in1                => s_in1(12,11),
			in2                => s_in2(12,11),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(11)
		);
	s_in1(12,11)            <= s_out1(13,11);
	s_in2(12,11)            <= s_out2(13,12);
	s_locks_lower_in(12,11) <= s_locks_lower_out(13,11);

		normal_cell_12_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,12),
			fetch              => s_fetch(12,12),
			data_in            => s_data_in(12,12),
			data_out           => s_data_out(12,12),
			out1               => s_out1(12,12),
			out2               => s_out2(12,12),
			lock_lower_row_out => s_locks_lower_out(12,12),
			lock_lower_row_in  => s_locks_lower_in(12,12),
			in1                => s_in1(12,12),
			in2                => s_in2(12,12),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(12)
		);
	s_in1(12,12)            <= s_out1(13,12);
	s_in2(12,12)            <= s_out2(13,13);
	s_locks_lower_in(12,12) <= s_locks_lower_out(13,12);

		normal_cell_12_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,13),
			fetch              => s_fetch(12,13),
			data_in            => s_data_in(12,13),
			data_out           => s_data_out(12,13),
			out1               => s_out1(12,13),
			out2               => s_out2(12,13),
			lock_lower_row_out => s_locks_lower_out(12,13),
			lock_lower_row_in  => s_locks_lower_in(12,13),
			in1                => s_in1(12,13),
			in2                => s_in2(12,13),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(13)
		);
	s_in1(12,13)            <= s_out1(13,13);
	s_in2(12,13)            <= s_out2(13,14);
	s_locks_lower_in(12,13) <= s_locks_lower_out(13,13);

		normal_cell_12_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,14),
			fetch              => s_fetch(12,14),
			data_in            => s_data_in(12,14),
			data_out           => s_data_out(12,14),
			out1               => s_out1(12,14),
			out2               => s_out2(12,14),
			lock_lower_row_out => s_locks_lower_out(12,14),
			lock_lower_row_in  => s_locks_lower_in(12,14),
			in1                => s_in1(12,14),
			in2                => s_in2(12,14),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(14)
		);
	s_in1(12,14)            <= s_out1(13,14);
	s_in2(12,14)            <= s_out2(13,15);
	s_locks_lower_in(12,14) <= s_locks_lower_out(13,14);

		normal_cell_12_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,15),
			fetch              => s_fetch(12,15),
			data_in            => s_data_in(12,15),
			data_out           => s_data_out(12,15),
			out1               => s_out1(12,15),
			out2               => s_out2(12,15),
			lock_lower_row_out => s_locks_lower_out(12,15),
			lock_lower_row_in  => s_locks_lower_in(12,15),
			in1                => s_in1(12,15),
			in2                => s_in2(12,15),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(15)
		);
	s_in1(12,15)            <= s_out1(13,15);
	s_in2(12,15)            <= s_out2(13,16);
	s_locks_lower_in(12,15) <= s_locks_lower_out(13,15);

		normal_cell_12_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,16),
			fetch              => s_fetch(12,16),
			data_in            => s_data_in(12,16),
			data_out           => s_data_out(12,16),
			out1               => s_out1(12,16),
			out2               => s_out2(12,16),
			lock_lower_row_out => s_locks_lower_out(12,16),
			lock_lower_row_in  => s_locks_lower_in(12,16),
			in1                => s_in1(12,16),
			in2                => s_in2(12,16),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(16)
		);
	s_in1(12,16)            <= s_out1(13,16);
	s_in2(12,16)            <= s_out2(13,17);
	s_locks_lower_in(12,16) <= s_locks_lower_out(13,16);

		normal_cell_12_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,17),
			fetch              => s_fetch(12,17),
			data_in            => s_data_in(12,17),
			data_out           => s_data_out(12,17),
			out1               => s_out1(12,17),
			out2               => s_out2(12,17),
			lock_lower_row_out => s_locks_lower_out(12,17),
			lock_lower_row_in  => s_locks_lower_in(12,17),
			in1                => s_in1(12,17),
			in2                => s_in2(12,17),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(17)
		);
	s_in1(12,17)            <= s_out1(13,17);
	s_in2(12,17)            <= s_out2(13,18);
	s_locks_lower_in(12,17) <= s_locks_lower_out(13,17);

		normal_cell_12_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,18),
			fetch              => s_fetch(12,18),
			data_in            => s_data_in(12,18),
			data_out           => s_data_out(12,18),
			out1               => s_out1(12,18),
			out2               => s_out2(12,18),
			lock_lower_row_out => s_locks_lower_out(12,18),
			lock_lower_row_in  => s_locks_lower_in(12,18),
			in1                => s_in1(12,18),
			in2                => s_in2(12,18),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(18)
		);
	s_in1(12,18)            <= s_out1(13,18);
	s_in2(12,18)            <= s_out2(13,19);
	s_locks_lower_in(12,18) <= s_locks_lower_out(13,18);

		normal_cell_12_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,19),
			fetch              => s_fetch(12,19),
			data_in            => s_data_in(12,19),
			data_out           => s_data_out(12,19),
			out1               => s_out1(12,19),
			out2               => s_out2(12,19),
			lock_lower_row_out => s_locks_lower_out(12,19),
			lock_lower_row_in  => s_locks_lower_in(12,19),
			in1                => s_in1(12,19),
			in2                => s_in2(12,19),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(19)
		);
	s_in1(12,19)            <= s_out1(13,19);
	s_in2(12,19)            <= s_out2(13,20);
	s_locks_lower_in(12,19) <= s_locks_lower_out(13,19);

		normal_cell_12_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,20),
			fetch              => s_fetch(12,20),
			data_in            => s_data_in(12,20),
			data_out           => s_data_out(12,20),
			out1               => s_out1(12,20),
			out2               => s_out2(12,20),
			lock_lower_row_out => s_locks_lower_out(12,20),
			lock_lower_row_in  => s_locks_lower_in(12,20),
			in1                => s_in1(12,20),
			in2                => s_in2(12,20),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(20)
		);
	s_in1(12,20)            <= s_out1(13,20);
	s_in2(12,20)            <= s_out2(13,21);
	s_locks_lower_in(12,20) <= s_locks_lower_out(13,20);

		normal_cell_12_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,21),
			fetch              => s_fetch(12,21),
			data_in            => s_data_in(12,21),
			data_out           => s_data_out(12,21),
			out1               => s_out1(12,21),
			out2               => s_out2(12,21),
			lock_lower_row_out => s_locks_lower_out(12,21),
			lock_lower_row_in  => s_locks_lower_in(12,21),
			in1                => s_in1(12,21),
			in2                => s_in2(12,21),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(21)
		);
	s_in1(12,21)            <= s_out1(13,21);
	s_in2(12,21)            <= s_out2(13,22);
	s_locks_lower_in(12,21) <= s_locks_lower_out(13,21);

		normal_cell_12_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,22),
			fetch              => s_fetch(12,22),
			data_in            => s_data_in(12,22),
			data_out           => s_data_out(12,22),
			out1               => s_out1(12,22),
			out2               => s_out2(12,22),
			lock_lower_row_out => s_locks_lower_out(12,22),
			lock_lower_row_in  => s_locks_lower_in(12,22),
			in1                => s_in1(12,22),
			in2                => s_in2(12,22),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(22)
		);
	s_in1(12,22)            <= s_out1(13,22);
	s_in2(12,22)            <= s_out2(13,23);
	s_locks_lower_in(12,22) <= s_locks_lower_out(13,22);

		normal_cell_12_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,23),
			fetch              => s_fetch(12,23),
			data_in            => s_data_in(12,23),
			data_out           => s_data_out(12,23),
			out1               => s_out1(12,23),
			out2               => s_out2(12,23),
			lock_lower_row_out => s_locks_lower_out(12,23),
			lock_lower_row_in  => s_locks_lower_in(12,23),
			in1                => s_in1(12,23),
			in2                => s_in2(12,23),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(23)
		);
	s_in1(12,23)            <= s_out1(13,23);
	s_in2(12,23)            <= s_out2(13,24);
	s_locks_lower_in(12,23) <= s_locks_lower_out(13,23);

		normal_cell_12_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,24),
			fetch              => s_fetch(12,24),
			data_in            => s_data_in(12,24),
			data_out           => s_data_out(12,24),
			out1               => s_out1(12,24),
			out2               => s_out2(12,24),
			lock_lower_row_out => s_locks_lower_out(12,24),
			lock_lower_row_in  => s_locks_lower_in(12,24),
			in1                => s_in1(12,24),
			in2                => s_in2(12,24),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(24)
		);
	s_in1(12,24)            <= s_out1(13,24);
	s_in2(12,24)            <= s_out2(13,25);
	s_locks_lower_in(12,24) <= s_locks_lower_out(13,24);

		normal_cell_12_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,25),
			fetch              => s_fetch(12,25),
			data_in            => s_data_in(12,25),
			data_out           => s_data_out(12,25),
			out1               => s_out1(12,25),
			out2               => s_out2(12,25),
			lock_lower_row_out => s_locks_lower_out(12,25),
			lock_lower_row_in  => s_locks_lower_in(12,25),
			in1                => s_in1(12,25),
			in2                => s_in2(12,25),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(25)
		);
	s_in1(12,25)            <= s_out1(13,25);
	s_in2(12,25)            <= s_out2(13,26);
	s_locks_lower_in(12,25) <= s_locks_lower_out(13,25);

		normal_cell_12_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,26),
			fetch              => s_fetch(12,26),
			data_in            => s_data_in(12,26),
			data_out           => s_data_out(12,26),
			out1               => s_out1(12,26),
			out2               => s_out2(12,26),
			lock_lower_row_out => s_locks_lower_out(12,26),
			lock_lower_row_in  => s_locks_lower_in(12,26),
			in1                => s_in1(12,26),
			in2                => s_in2(12,26),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(26)
		);
	s_in1(12,26)            <= s_out1(13,26);
	s_in2(12,26)            <= s_out2(13,27);
	s_locks_lower_in(12,26) <= s_locks_lower_out(13,26);

		normal_cell_12_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,27),
			fetch              => s_fetch(12,27),
			data_in            => s_data_in(12,27),
			data_out           => s_data_out(12,27),
			out1               => s_out1(12,27),
			out2               => s_out2(12,27),
			lock_lower_row_out => s_locks_lower_out(12,27),
			lock_lower_row_in  => s_locks_lower_in(12,27),
			in1                => s_in1(12,27),
			in2                => s_in2(12,27),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(27)
		);
	s_in1(12,27)            <= s_out1(13,27);
	s_in2(12,27)            <= s_out2(13,28);
	s_locks_lower_in(12,27) <= s_locks_lower_out(13,27);

		normal_cell_12_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,28),
			fetch              => s_fetch(12,28),
			data_in            => s_data_in(12,28),
			data_out           => s_data_out(12,28),
			out1               => s_out1(12,28),
			out2               => s_out2(12,28),
			lock_lower_row_out => s_locks_lower_out(12,28),
			lock_lower_row_in  => s_locks_lower_in(12,28),
			in1                => s_in1(12,28),
			in2                => s_in2(12,28),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(28)
		);
	s_in1(12,28)            <= s_out1(13,28);
	s_in2(12,28)            <= s_out2(13,29);
	s_locks_lower_in(12,28) <= s_locks_lower_out(13,28);

		normal_cell_12_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,29),
			fetch              => s_fetch(12,29),
			data_in            => s_data_in(12,29),
			data_out           => s_data_out(12,29),
			out1               => s_out1(12,29),
			out2               => s_out2(12,29),
			lock_lower_row_out => s_locks_lower_out(12,29),
			lock_lower_row_in  => s_locks_lower_in(12,29),
			in1                => s_in1(12,29),
			in2                => s_in2(12,29),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(29)
		);
	s_in1(12,29)            <= s_out1(13,29);
	s_in2(12,29)            <= s_out2(13,30);
	s_locks_lower_in(12,29) <= s_locks_lower_out(13,29);

		normal_cell_12_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,30),
			fetch              => s_fetch(12,30),
			data_in            => s_data_in(12,30),
			data_out           => s_data_out(12,30),
			out1               => s_out1(12,30),
			out2               => s_out2(12,30),
			lock_lower_row_out => s_locks_lower_out(12,30),
			lock_lower_row_in  => s_locks_lower_in(12,30),
			in1                => s_in1(12,30),
			in2                => s_in2(12,30),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(30)
		);
	s_in1(12,30)            <= s_out1(13,30);
	s_in2(12,30)            <= s_out2(13,31);
	s_locks_lower_in(12,30) <= s_locks_lower_out(13,30);

		normal_cell_12_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,31),
			fetch              => s_fetch(12,31),
			data_in            => s_data_in(12,31),
			data_out           => s_data_out(12,31),
			out1               => s_out1(12,31),
			out2               => s_out2(12,31),
			lock_lower_row_out => s_locks_lower_out(12,31),
			lock_lower_row_in  => s_locks_lower_in(12,31),
			in1                => s_in1(12,31),
			in2                => s_in2(12,31),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(31)
		);
	s_in1(12,31)            <= s_out1(13,31);
	s_in2(12,31)            <= s_out2(13,32);
	s_locks_lower_in(12,31) <= s_locks_lower_out(13,31);

		normal_cell_12_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,32),
			fetch              => s_fetch(12,32),
			data_in            => s_data_in(12,32),
			data_out           => s_data_out(12,32),
			out1               => s_out1(12,32),
			out2               => s_out2(12,32),
			lock_lower_row_out => s_locks_lower_out(12,32),
			lock_lower_row_in  => s_locks_lower_in(12,32),
			in1                => s_in1(12,32),
			in2                => s_in2(12,32),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(32)
		);
	s_in1(12,32)            <= s_out1(13,32);
	s_in2(12,32)            <= s_out2(13,33);
	s_locks_lower_in(12,32) <= s_locks_lower_out(13,32);

		normal_cell_12_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,33),
			fetch              => s_fetch(12,33),
			data_in            => s_data_in(12,33),
			data_out           => s_data_out(12,33),
			out1               => s_out1(12,33),
			out2               => s_out2(12,33),
			lock_lower_row_out => s_locks_lower_out(12,33),
			lock_lower_row_in  => s_locks_lower_in(12,33),
			in1                => s_in1(12,33),
			in2                => s_in2(12,33),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(33)
		);
	s_in1(12,33)            <= s_out1(13,33);
	s_in2(12,33)            <= s_out2(13,34);
	s_locks_lower_in(12,33) <= s_locks_lower_out(13,33);

		normal_cell_12_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,34),
			fetch              => s_fetch(12,34),
			data_in            => s_data_in(12,34),
			data_out           => s_data_out(12,34),
			out1               => s_out1(12,34),
			out2               => s_out2(12,34),
			lock_lower_row_out => s_locks_lower_out(12,34),
			lock_lower_row_in  => s_locks_lower_in(12,34),
			in1                => s_in1(12,34),
			in2                => s_in2(12,34),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(34)
		);
	s_in1(12,34)            <= s_out1(13,34);
	s_in2(12,34)            <= s_out2(13,35);
	s_locks_lower_in(12,34) <= s_locks_lower_out(13,34);

		normal_cell_12_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,35),
			fetch              => s_fetch(12,35),
			data_in            => s_data_in(12,35),
			data_out           => s_data_out(12,35),
			out1               => s_out1(12,35),
			out2               => s_out2(12,35),
			lock_lower_row_out => s_locks_lower_out(12,35),
			lock_lower_row_in  => s_locks_lower_in(12,35),
			in1                => s_in1(12,35),
			in2                => s_in2(12,35),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(35)
		);
	s_in1(12,35)            <= s_out1(13,35);
	s_in2(12,35)            <= s_out2(13,36);
	s_locks_lower_in(12,35) <= s_locks_lower_out(13,35);

		normal_cell_12_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,36),
			fetch              => s_fetch(12,36),
			data_in            => s_data_in(12,36),
			data_out           => s_data_out(12,36),
			out1               => s_out1(12,36),
			out2               => s_out2(12,36),
			lock_lower_row_out => s_locks_lower_out(12,36),
			lock_lower_row_in  => s_locks_lower_in(12,36),
			in1                => s_in1(12,36),
			in2                => s_in2(12,36),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(36)
		);
	s_in1(12,36)            <= s_out1(13,36);
	s_in2(12,36)            <= s_out2(13,37);
	s_locks_lower_in(12,36) <= s_locks_lower_out(13,36);

		normal_cell_12_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,37),
			fetch              => s_fetch(12,37),
			data_in            => s_data_in(12,37),
			data_out           => s_data_out(12,37),
			out1               => s_out1(12,37),
			out2               => s_out2(12,37),
			lock_lower_row_out => s_locks_lower_out(12,37),
			lock_lower_row_in  => s_locks_lower_in(12,37),
			in1                => s_in1(12,37),
			in2                => s_in2(12,37),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(37)
		);
	s_in1(12,37)            <= s_out1(13,37);
	s_in2(12,37)            <= s_out2(13,38);
	s_locks_lower_in(12,37) <= s_locks_lower_out(13,37);

		normal_cell_12_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,38),
			fetch              => s_fetch(12,38),
			data_in            => s_data_in(12,38),
			data_out           => s_data_out(12,38),
			out1               => s_out1(12,38),
			out2               => s_out2(12,38),
			lock_lower_row_out => s_locks_lower_out(12,38),
			lock_lower_row_in  => s_locks_lower_in(12,38),
			in1                => s_in1(12,38),
			in2                => s_in2(12,38),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(38)
		);
	s_in1(12,38)            <= s_out1(13,38);
	s_in2(12,38)            <= s_out2(13,39);
	s_locks_lower_in(12,38) <= s_locks_lower_out(13,38);

		normal_cell_12_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,39),
			fetch              => s_fetch(12,39),
			data_in            => s_data_in(12,39),
			data_out           => s_data_out(12,39),
			out1               => s_out1(12,39),
			out2               => s_out2(12,39),
			lock_lower_row_out => s_locks_lower_out(12,39),
			lock_lower_row_in  => s_locks_lower_in(12,39),
			in1                => s_in1(12,39),
			in2                => s_in2(12,39),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(39)
		);
	s_in1(12,39)            <= s_out1(13,39);
	s_in2(12,39)            <= s_out2(13,40);
	s_locks_lower_in(12,39) <= s_locks_lower_out(13,39);

		normal_cell_12_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,40),
			fetch              => s_fetch(12,40),
			data_in            => s_data_in(12,40),
			data_out           => s_data_out(12,40),
			out1               => s_out1(12,40),
			out2               => s_out2(12,40),
			lock_lower_row_out => s_locks_lower_out(12,40),
			lock_lower_row_in  => s_locks_lower_in(12,40),
			in1                => s_in1(12,40),
			in2                => s_in2(12,40),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(40)
		);
	s_in1(12,40)            <= s_out1(13,40);
	s_in2(12,40)            <= s_out2(13,41);
	s_locks_lower_in(12,40) <= s_locks_lower_out(13,40);

		normal_cell_12_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,41),
			fetch              => s_fetch(12,41),
			data_in            => s_data_in(12,41),
			data_out           => s_data_out(12,41),
			out1               => s_out1(12,41),
			out2               => s_out2(12,41),
			lock_lower_row_out => s_locks_lower_out(12,41),
			lock_lower_row_in  => s_locks_lower_in(12,41),
			in1                => s_in1(12,41),
			in2                => s_in2(12,41),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(41)
		);
	s_in1(12,41)            <= s_out1(13,41);
	s_in2(12,41)            <= s_out2(13,42);
	s_locks_lower_in(12,41) <= s_locks_lower_out(13,41);

		normal_cell_12_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,42),
			fetch              => s_fetch(12,42),
			data_in            => s_data_in(12,42),
			data_out           => s_data_out(12,42),
			out1               => s_out1(12,42),
			out2               => s_out2(12,42),
			lock_lower_row_out => s_locks_lower_out(12,42),
			lock_lower_row_in  => s_locks_lower_in(12,42),
			in1                => s_in1(12,42),
			in2                => s_in2(12,42),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(42)
		);
	s_in1(12,42)            <= s_out1(13,42);
	s_in2(12,42)            <= s_out2(13,43);
	s_locks_lower_in(12,42) <= s_locks_lower_out(13,42);

		normal_cell_12_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,43),
			fetch              => s_fetch(12,43),
			data_in            => s_data_in(12,43),
			data_out           => s_data_out(12,43),
			out1               => s_out1(12,43),
			out2               => s_out2(12,43),
			lock_lower_row_out => s_locks_lower_out(12,43),
			lock_lower_row_in  => s_locks_lower_in(12,43),
			in1                => s_in1(12,43),
			in2                => s_in2(12,43),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(43)
		);
	s_in1(12,43)            <= s_out1(13,43);
	s_in2(12,43)            <= s_out2(13,44);
	s_locks_lower_in(12,43) <= s_locks_lower_out(13,43);

		normal_cell_12_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,44),
			fetch              => s_fetch(12,44),
			data_in            => s_data_in(12,44),
			data_out           => s_data_out(12,44),
			out1               => s_out1(12,44),
			out2               => s_out2(12,44),
			lock_lower_row_out => s_locks_lower_out(12,44),
			lock_lower_row_in  => s_locks_lower_in(12,44),
			in1                => s_in1(12,44),
			in2                => s_in2(12,44),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(44)
		);
	s_in1(12,44)            <= s_out1(13,44);
	s_in2(12,44)            <= s_out2(13,45);
	s_locks_lower_in(12,44) <= s_locks_lower_out(13,44);

		normal_cell_12_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,45),
			fetch              => s_fetch(12,45),
			data_in            => s_data_in(12,45),
			data_out           => s_data_out(12,45),
			out1               => s_out1(12,45),
			out2               => s_out2(12,45),
			lock_lower_row_out => s_locks_lower_out(12,45),
			lock_lower_row_in  => s_locks_lower_in(12,45),
			in1                => s_in1(12,45),
			in2                => s_in2(12,45),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(45)
		);
	s_in1(12,45)            <= s_out1(13,45);
	s_in2(12,45)            <= s_out2(13,46);
	s_locks_lower_in(12,45) <= s_locks_lower_out(13,45);

		normal_cell_12_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,46),
			fetch              => s_fetch(12,46),
			data_in            => s_data_in(12,46),
			data_out           => s_data_out(12,46),
			out1               => s_out1(12,46),
			out2               => s_out2(12,46),
			lock_lower_row_out => s_locks_lower_out(12,46),
			lock_lower_row_in  => s_locks_lower_in(12,46),
			in1                => s_in1(12,46),
			in2                => s_in2(12,46),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(46)
		);
	s_in1(12,46)            <= s_out1(13,46);
	s_in2(12,46)            <= s_out2(13,47);
	s_locks_lower_in(12,46) <= s_locks_lower_out(13,46);

		normal_cell_12_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,47),
			fetch              => s_fetch(12,47),
			data_in            => s_data_in(12,47),
			data_out           => s_data_out(12,47),
			out1               => s_out1(12,47),
			out2               => s_out2(12,47),
			lock_lower_row_out => s_locks_lower_out(12,47),
			lock_lower_row_in  => s_locks_lower_in(12,47),
			in1                => s_in1(12,47),
			in2                => s_in2(12,47),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(47)
		);
	s_in1(12,47)            <= s_out1(13,47);
	s_in2(12,47)            <= s_out2(13,48);
	s_locks_lower_in(12,47) <= s_locks_lower_out(13,47);

		normal_cell_12_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,48),
			fetch              => s_fetch(12,48),
			data_in            => s_data_in(12,48),
			data_out           => s_data_out(12,48),
			out1               => s_out1(12,48),
			out2               => s_out2(12,48),
			lock_lower_row_out => s_locks_lower_out(12,48),
			lock_lower_row_in  => s_locks_lower_in(12,48),
			in1                => s_in1(12,48),
			in2                => s_in2(12,48),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(48)
		);
	s_in1(12,48)            <= s_out1(13,48);
	s_in2(12,48)            <= s_out2(13,49);
	s_locks_lower_in(12,48) <= s_locks_lower_out(13,48);

		normal_cell_12_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,49),
			fetch              => s_fetch(12,49),
			data_in            => s_data_in(12,49),
			data_out           => s_data_out(12,49),
			out1               => s_out1(12,49),
			out2               => s_out2(12,49),
			lock_lower_row_out => s_locks_lower_out(12,49),
			lock_lower_row_in  => s_locks_lower_in(12,49),
			in1                => s_in1(12,49),
			in2                => s_in2(12,49),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(49)
		);
	s_in1(12,49)            <= s_out1(13,49);
	s_in2(12,49)            <= s_out2(13,50);
	s_locks_lower_in(12,49) <= s_locks_lower_out(13,49);

		normal_cell_12_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,50),
			fetch              => s_fetch(12,50),
			data_in            => s_data_in(12,50),
			data_out           => s_data_out(12,50),
			out1               => s_out1(12,50),
			out2               => s_out2(12,50),
			lock_lower_row_out => s_locks_lower_out(12,50),
			lock_lower_row_in  => s_locks_lower_in(12,50),
			in1                => s_in1(12,50),
			in2                => s_in2(12,50),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(50)
		);
	s_in1(12,50)            <= s_out1(13,50);
	s_in2(12,50)            <= s_out2(13,51);
	s_locks_lower_in(12,50) <= s_locks_lower_out(13,50);

		normal_cell_12_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,51),
			fetch              => s_fetch(12,51),
			data_in            => s_data_in(12,51),
			data_out           => s_data_out(12,51),
			out1               => s_out1(12,51),
			out2               => s_out2(12,51),
			lock_lower_row_out => s_locks_lower_out(12,51),
			lock_lower_row_in  => s_locks_lower_in(12,51),
			in1                => s_in1(12,51),
			in2                => s_in2(12,51),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(51)
		);
	s_in1(12,51)            <= s_out1(13,51);
	s_in2(12,51)            <= s_out2(13,52);
	s_locks_lower_in(12,51) <= s_locks_lower_out(13,51);

		normal_cell_12_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,52),
			fetch              => s_fetch(12,52),
			data_in            => s_data_in(12,52),
			data_out           => s_data_out(12,52),
			out1               => s_out1(12,52),
			out2               => s_out2(12,52),
			lock_lower_row_out => s_locks_lower_out(12,52),
			lock_lower_row_in  => s_locks_lower_in(12,52),
			in1                => s_in1(12,52),
			in2                => s_in2(12,52),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(52)
		);
	s_in1(12,52)            <= s_out1(13,52);
	s_in2(12,52)            <= s_out2(13,53);
	s_locks_lower_in(12,52) <= s_locks_lower_out(13,52);

		normal_cell_12_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,53),
			fetch              => s_fetch(12,53),
			data_in            => s_data_in(12,53),
			data_out           => s_data_out(12,53),
			out1               => s_out1(12,53),
			out2               => s_out2(12,53),
			lock_lower_row_out => s_locks_lower_out(12,53),
			lock_lower_row_in  => s_locks_lower_in(12,53),
			in1                => s_in1(12,53),
			in2                => s_in2(12,53),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(53)
		);
	s_in1(12,53)            <= s_out1(13,53);
	s_in2(12,53)            <= s_out2(13,54);
	s_locks_lower_in(12,53) <= s_locks_lower_out(13,53);

		normal_cell_12_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,54),
			fetch              => s_fetch(12,54),
			data_in            => s_data_in(12,54),
			data_out           => s_data_out(12,54),
			out1               => s_out1(12,54),
			out2               => s_out2(12,54),
			lock_lower_row_out => s_locks_lower_out(12,54),
			lock_lower_row_in  => s_locks_lower_in(12,54),
			in1                => s_in1(12,54),
			in2                => s_in2(12,54),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(54)
		);
	s_in1(12,54)            <= s_out1(13,54);
	s_in2(12,54)            <= s_out2(13,55);
	s_locks_lower_in(12,54) <= s_locks_lower_out(13,54);

		normal_cell_12_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,55),
			fetch              => s_fetch(12,55),
			data_in            => s_data_in(12,55),
			data_out           => s_data_out(12,55),
			out1               => s_out1(12,55),
			out2               => s_out2(12,55),
			lock_lower_row_out => s_locks_lower_out(12,55),
			lock_lower_row_in  => s_locks_lower_in(12,55),
			in1                => s_in1(12,55),
			in2                => s_in2(12,55),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(55)
		);
	s_in1(12,55)            <= s_out1(13,55);
	s_in2(12,55)            <= s_out2(13,56);
	s_locks_lower_in(12,55) <= s_locks_lower_out(13,55);

		normal_cell_12_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,56),
			fetch              => s_fetch(12,56),
			data_in            => s_data_in(12,56),
			data_out           => s_data_out(12,56),
			out1               => s_out1(12,56),
			out2               => s_out2(12,56),
			lock_lower_row_out => s_locks_lower_out(12,56),
			lock_lower_row_in  => s_locks_lower_in(12,56),
			in1                => s_in1(12,56),
			in2                => s_in2(12,56),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(56)
		);
	s_in1(12,56)            <= s_out1(13,56);
	s_in2(12,56)            <= s_out2(13,57);
	s_locks_lower_in(12,56) <= s_locks_lower_out(13,56);

		normal_cell_12_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,57),
			fetch              => s_fetch(12,57),
			data_in            => s_data_in(12,57),
			data_out           => s_data_out(12,57),
			out1               => s_out1(12,57),
			out2               => s_out2(12,57),
			lock_lower_row_out => s_locks_lower_out(12,57),
			lock_lower_row_in  => s_locks_lower_in(12,57),
			in1                => s_in1(12,57),
			in2                => s_in2(12,57),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(57)
		);
	s_in1(12,57)            <= s_out1(13,57);
	s_in2(12,57)            <= s_out2(13,58);
	s_locks_lower_in(12,57) <= s_locks_lower_out(13,57);

		normal_cell_12_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,58),
			fetch              => s_fetch(12,58),
			data_in            => s_data_in(12,58),
			data_out           => s_data_out(12,58),
			out1               => s_out1(12,58),
			out2               => s_out2(12,58),
			lock_lower_row_out => s_locks_lower_out(12,58),
			lock_lower_row_in  => s_locks_lower_in(12,58),
			in1                => s_in1(12,58),
			in2                => s_in2(12,58),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(58)
		);
	s_in1(12,58)            <= s_out1(13,58);
	s_in2(12,58)            <= s_out2(13,59);
	s_locks_lower_in(12,58) <= s_locks_lower_out(13,58);

		normal_cell_12_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,59),
			fetch              => s_fetch(12,59),
			data_in            => s_data_in(12,59),
			data_out           => s_data_out(12,59),
			out1               => s_out1(12,59),
			out2               => s_out2(12,59),
			lock_lower_row_out => s_locks_lower_out(12,59),
			lock_lower_row_in  => s_locks_lower_in(12,59),
			in1                => s_in1(12,59),
			in2                => s_in2(12,59),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(59)
		);
	s_in1(12,59)            <= s_out1(13,59);
	s_in2(12,59)            <= s_out2(13,60);
	s_locks_lower_in(12,59) <= s_locks_lower_out(13,59);

		last_col_cell_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(12,60),
			fetch              => s_fetch(12,60),
			data_in            => s_data_in(12,60),
			data_out           => s_data_out(12,60),
			out1               => s_out1(12,60),
			out2               => s_out2(12,60),
			lock_lower_row_out => s_locks_lower_out(12,60),
			lock_lower_row_in  => s_locks_lower_in(12,60),
			in1                => s_in1(12,60),
			in2                => (others => '0'),
			lock_row           => s_locks(12),
			piv_found          => s_piv_found,
			row_data           => s_row_data(12),
			col_data           => s_col_data(60)
		);
	s_in1(12,60)            <= s_out1(13,60);
	s_locks_lower_in(12,60) <= s_locks_lower_out(13,60);

		normal_cell_13_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,1),
			fetch              => s_fetch(13,1),
			data_in            => s_data_in(13,1),
			data_out           => s_data_out(13,1),
			out1               => s_out1(13,1),
			out2               => s_out2(13,1),
			lock_lower_row_out => s_locks_lower_out(13,1),
			lock_lower_row_in  => s_locks_lower_in(13,1),
			in1                => s_in1(13,1),
			in2                => s_in2(13,1),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(1)
		);
	s_in1(13,1)            <= s_out1(14,1);
	s_in2(13,1)            <= s_out2(14,2);
	s_locks_lower_in(13,1) <= s_locks_lower_out(14,1);

		normal_cell_13_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,2),
			fetch              => s_fetch(13,2),
			data_in            => s_data_in(13,2),
			data_out           => s_data_out(13,2),
			out1               => s_out1(13,2),
			out2               => s_out2(13,2),
			lock_lower_row_out => s_locks_lower_out(13,2),
			lock_lower_row_in  => s_locks_lower_in(13,2),
			in1                => s_in1(13,2),
			in2                => s_in2(13,2),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(2)
		);
	s_in1(13,2)            <= s_out1(14,2);
	s_in2(13,2)            <= s_out2(14,3);
	s_locks_lower_in(13,2) <= s_locks_lower_out(14,2);

		normal_cell_13_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,3),
			fetch              => s_fetch(13,3),
			data_in            => s_data_in(13,3),
			data_out           => s_data_out(13,3),
			out1               => s_out1(13,3),
			out2               => s_out2(13,3),
			lock_lower_row_out => s_locks_lower_out(13,3),
			lock_lower_row_in  => s_locks_lower_in(13,3),
			in1                => s_in1(13,3),
			in2                => s_in2(13,3),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(3)
		);
	s_in1(13,3)            <= s_out1(14,3);
	s_in2(13,3)            <= s_out2(14,4);
	s_locks_lower_in(13,3) <= s_locks_lower_out(14,3);

		normal_cell_13_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,4),
			fetch              => s_fetch(13,4),
			data_in            => s_data_in(13,4),
			data_out           => s_data_out(13,4),
			out1               => s_out1(13,4),
			out2               => s_out2(13,4),
			lock_lower_row_out => s_locks_lower_out(13,4),
			lock_lower_row_in  => s_locks_lower_in(13,4),
			in1                => s_in1(13,4),
			in2                => s_in2(13,4),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(4)
		);
	s_in1(13,4)            <= s_out1(14,4);
	s_in2(13,4)            <= s_out2(14,5);
	s_locks_lower_in(13,4) <= s_locks_lower_out(14,4);

		normal_cell_13_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,5),
			fetch              => s_fetch(13,5),
			data_in            => s_data_in(13,5),
			data_out           => s_data_out(13,5),
			out1               => s_out1(13,5),
			out2               => s_out2(13,5),
			lock_lower_row_out => s_locks_lower_out(13,5),
			lock_lower_row_in  => s_locks_lower_in(13,5),
			in1                => s_in1(13,5),
			in2                => s_in2(13,5),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(5)
		);
	s_in1(13,5)            <= s_out1(14,5);
	s_in2(13,5)            <= s_out2(14,6);
	s_locks_lower_in(13,5) <= s_locks_lower_out(14,5);

		normal_cell_13_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,6),
			fetch              => s_fetch(13,6),
			data_in            => s_data_in(13,6),
			data_out           => s_data_out(13,6),
			out1               => s_out1(13,6),
			out2               => s_out2(13,6),
			lock_lower_row_out => s_locks_lower_out(13,6),
			lock_lower_row_in  => s_locks_lower_in(13,6),
			in1                => s_in1(13,6),
			in2                => s_in2(13,6),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(6)
		);
	s_in1(13,6)            <= s_out1(14,6);
	s_in2(13,6)            <= s_out2(14,7);
	s_locks_lower_in(13,6) <= s_locks_lower_out(14,6);

		normal_cell_13_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,7),
			fetch              => s_fetch(13,7),
			data_in            => s_data_in(13,7),
			data_out           => s_data_out(13,7),
			out1               => s_out1(13,7),
			out2               => s_out2(13,7),
			lock_lower_row_out => s_locks_lower_out(13,7),
			lock_lower_row_in  => s_locks_lower_in(13,7),
			in1                => s_in1(13,7),
			in2                => s_in2(13,7),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(7)
		);
	s_in1(13,7)            <= s_out1(14,7);
	s_in2(13,7)            <= s_out2(14,8);
	s_locks_lower_in(13,7) <= s_locks_lower_out(14,7);

		normal_cell_13_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,8),
			fetch              => s_fetch(13,8),
			data_in            => s_data_in(13,8),
			data_out           => s_data_out(13,8),
			out1               => s_out1(13,8),
			out2               => s_out2(13,8),
			lock_lower_row_out => s_locks_lower_out(13,8),
			lock_lower_row_in  => s_locks_lower_in(13,8),
			in1                => s_in1(13,8),
			in2                => s_in2(13,8),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(8)
		);
	s_in1(13,8)            <= s_out1(14,8);
	s_in2(13,8)            <= s_out2(14,9);
	s_locks_lower_in(13,8) <= s_locks_lower_out(14,8);

		normal_cell_13_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,9),
			fetch              => s_fetch(13,9),
			data_in            => s_data_in(13,9),
			data_out           => s_data_out(13,9),
			out1               => s_out1(13,9),
			out2               => s_out2(13,9),
			lock_lower_row_out => s_locks_lower_out(13,9),
			lock_lower_row_in  => s_locks_lower_in(13,9),
			in1                => s_in1(13,9),
			in2                => s_in2(13,9),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(9)
		);
	s_in1(13,9)            <= s_out1(14,9);
	s_in2(13,9)            <= s_out2(14,10);
	s_locks_lower_in(13,9) <= s_locks_lower_out(14,9);

		normal_cell_13_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,10),
			fetch              => s_fetch(13,10),
			data_in            => s_data_in(13,10),
			data_out           => s_data_out(13,10),
			out1               => s_out1(13,10),
			out2               => s_out2(13,10),
			lock_lower_row_out => s_locks_lower_out(13,10),
			lock_lower_row_in  => s_locks_lower_in(13,10),
			in1                => s_in1(13,10),
			in2                => s_in2(13,10),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(10)
		);
	s_in1(13,10)            <= s_out1(14,10);
	s_in2(13,10)            <= s_out2(14,11);
	s_locks_lower_in(13,10) <= s_locks_lower_out(14,10);

		normal_cell_13_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,11),
			fetch              => s_fetch(13,11),
			data_in            => s_data_in(13,11),
			data_out           => s_data_out(13,11),
			out1               => s_out1(13,11),
			out2               => s_out2(13,11),
			lock_lower_row_out => s_locks_lower_out(13,11),
			lock_lower_row_in  => s_locks_lower_in(13,11),
			in1                => s_in1(13,11),
			in2                => s_in2(13,11),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(11)
		);
	s_in1(13,11)            <= s_out1(14,11);
	s_in2(13,11)            <= s_out2(14,12);
	s_locks_lower_in(13,11) <= s_locks_lower_out(14,11);

		normal_cell_13_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,12),
			fetch              => s_fetch(13,12),
			data_in            => s_data_in(13,12),
			data_out           => s_data_out(13,12),
			out1               => s_out1(13,12),
			out2               => s_out2(13,12),
			lock_lower_row_out => s_locks_lower_out(13,12),
			lock_lower_row_in  => s_locks_lower_in(13,12),
			in1                => s_in1(13,12),
			in2                => s_in2(13,12),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(12)
		);
	s_in1(13,12)            <= s_out1(14,12);
	s_in2(13,12)            <= s_out2(14,13);
	s_locks_lower_in(13,12) <= s_locks_lower_out(14,12);

		normal_cell_13_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,13),
			fetch              => s_fetch(13,13),
			data_in            => s_data_in(13,13),
			data_out           => s_data_out(13,13),
			out1               => s_out1(13,13),
			out2               => s_out2(13,13),
			lock_lower_row_out => s_locks_lower_out(13,13),
			lock_lower_row_in  => s_locks_lower_in(13,13),
			in1                => s_in1(13,13),
			in2                => s_in2(13,13),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(13)
		);
	s_in1(13,13)            <= s_out1(14,13);
	s_in2(13,13)            <= s_out2(14,14);
	s_locks_lower_in(13,13) <= s_locks_lower_out(14,13);

		normal_cell_13_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,14),
			fetch              => s_fetch(13,14),
			data_in            => s_data_in(13,14),
			data_out           => s_data_out(13,14),
			out1               => s_out1(13,14),
			out2               => s_out2(13,14),
			lock_lower_row_out => s_locks_lower_out(13,14),
			lock_lower_row_in  => s_locks_lower_in(13,14),
			in1                => s_in1(13,14),
			in2                => s_in2(13,14),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(14)
		);
	s_in1(13,14)            <= s_out1(14,14);
	s_in2(13,14)            <= s_out2(14,15);
	s_locks_lower_in(13,14) <= s_locks_lower_out(14,14);

		normal_cell_13_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,15),
			fetch              => s_fetch(13,15),
			data_in            => s_data_in(13,15),
			data_out           => s_data_out(13,15),
			out1               => s_out1(13,15),
			out2               => s_out2(13,15),
			lock_lower_row_out => s_locks_lower_out(13,15),
			lock_lower_row_in  => s_locks_lower_in(13,15),
			in1                => s_in1(13,15),
			in2                => s_in2(13,15),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(15)
		);
	s_in1(13,15)            <= s_out1(14,15);
	s_in2(13,15)            <= s_out2(14,16);
	s_locks_lower_in(13,15) <= s_locks_lower_out(14,15);

		normal_cell_13_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,16),
			fetch              => s_fetch(13,16),
			data_in            => s_data_in(13,16),
			data_out           => s_data_out(13,16),
			out1               => s_out1(13,16),
			out2               => s_out2(13,16),
			lock_lower_row_out => s_locks_lower_out(13,16),
			lock_lower_row_in  => s_locks_lower_in(13,16),
			in1                => s_in1(13,16),
			in2                => s_in2(13,16),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(16)
		);
	s_in1(13,16)            <= s_out1(14,16);
	s_in2(13,16)            <= s_out2(14,17);
	s_locks_lower_in(13,16) <= s_locks_lower_out(14,16);

		normal_cell_13_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,17),
			fetch              => s_fetch(13,17),
			data_in            => s_data_in(13,17),
			data_out           => s_data_out(13,17),
			out1               => s_out1(13,17),
			out2               => s_out2(13,17),
			lock_lower_row_out => s_locks_lower_out(13,17),
			lock_lower_row_in  => s_locks_lower_in(13,17),
			in1                => s_in1(13,17),
			in2                => s_in2(13,17),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(17)
		);
	s_in1(13,17)            <= s_out1(14,17);
	s_in2(13,17)            <= s_out2(14,18);
	s_locks_lower_in(13,17) <= s_locks_lower_out(14,17);

		normal_cell_13_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,18),
			fetch              => s_fetch(13,18),
			data_in            => s_data_in(13,18),
			data_out           => s_data_out(13,18),
			out1               => s_out1(13,18),
			out2               => s_out2(13,18),
			lock_lower_row_out => s_locks_lower_out(13,18),
			lock_lower_row_in  => s_locks_lower_in(13,18),
			in1                => s_in1(13,18),
			in2                => s_in2(13,18),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(18)
		);
	s_in1(13,18)            <= s_out1(14,18);
	s_in2(13,18)            <= s_out2(14,19);
	s_locks_lower_in(13,18) <= s_locks_lower_out(14,18);

		normal_cell_13_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,19),
			fetch              => s_fetch(13,19),
			data_in            => s_data_in(13,19),
			data_out           => s_data_out(13,19),
			out1               => s_out1(13,19),
			out2               => s_out2(13,19),
			lock_lower_row_out => s_locks_lower_out(13,19),
			lock_lower_row_in  => s_locks_lower_in(13,19),
			in1                => s_in1(13,19),
			in2                => s_in2(13,19),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(19)
		);
	s_in1(13,19)            <= s_out1(14,19);
	s_in2(13,19)            <= s_out2(14,20);
	s_locks_lower_in(13,19) <= s_locks_lower_out(14,19);

		normal_cell_13_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,20),
			fetch              => s_fetch(13,20),
			data_in            => s_data_in(13,20),
			data_out           => s_data_out(13,20),
			out1               => s_out1(13,20),
			out2               => s_out2(13,20),
			lock_lower_row_out => s_locks_lower_out(13,20),
			lock_lower_row_in  => s_locks_lower_in(13,20),
			in1                => s_in1(13,20),
			in2                => s_in2(13,20),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(20)
		);
	s_in1(13,20)            <= s_out1(14,20);
	s_in2(13,20)            <= s_out2(14,21);
	s_locks_lower_in(13,20) <= s_locks_lower_out(14,20);

		normal_cell_13_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,21),
			fetch              => s_fetch(13,21),
			data_in            => s_data_in(13,21),
			data_out           => s_data_out(13,21),
			out1               => s_out1(13,21),
			out2               => s_out2(13,21),
			lock_lower_row_out => s_locks_lower_out(13,21),
			lock_lower_row_in  => s_locks_lower_in(13,21),
			in1                => s_in1(13,21),
			in2                => s_in2(13,21),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(21)
		);
	s_in1(13,21)            <= s_out1(14,21);
	s_in2(13,21)            <= s_out2(14,22);
	s_locks_lower_in(13,21) <= s_locks_lower_out(14,21);

		normal_cell_13_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,22),
			fetch              => s_fetch(13,22),
			data_in            => s_data_in(13,22),
			data_out           => s_data_out(13,22),
			out1               => s_out1(13,22),
			out2               => s_out2(13,22),
			lock_lower_row_out => s_locks_lower_out(13,22),
			lock_lower_row_in  => s_locks_lower_in(13,22),
			in1                => s_in1(13,22),
			in2                => s_in2(13,22),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(22)
		);
	s_in1(13,22)            <= s_out1(14,22);
	s_in2(13,22)            <= s_out2(14,23);
	s_locks_lower_in(13,22) <= s_locks_lower_out(14,22);

		normal_cell_13_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,23),
			fetch              => s_fetch(13,23),
			data_in            => s_data_in(13,23),
			data_out           => s_data_out(13,23),
			out1               => s_out1(13,23),
			out2               => s_out2(13,23),
			lock_lower_row_out => s_locks_lower_out(13,23),
			lock_lower_row_in  => s_locks_lower_in(13,23),
			in1                => s_in1(13,23),
			in2                => s_in2(13,23),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(23)
		);
	s_in1(13,23)            <= s_out1(14,23);
	s_in2(13,23)            <= s_out2(14,24);
	s_locks_lower_in(13,23) <= s_locks_lower_out(14,23);

		normal_cell_13_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,24),
			fetch              => s_fetch(13,24),
			data_in            => s_data_in(13,24),
			data_out           => s_data_out(13,24),
			out1               => s_out1(13,24),
			out2               => s_out2(13,24),
			lock_lower_row_out => s_locks_lower_out(13,24),
			lock_lower_row_in  => s_locks_lower_in(13,24),
			in1                => s_in1(13,24),
			in2                => s_in2(13,24),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(24)
		);
	s_in1(13,24)            <= s_out1(14,24);
	s_in2(13,24)            <= s_out2(14,25);
	s_locks_lower_in(13,24) <= s_locks_lower_out(14,24);

		normal_cell_13_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,25),
			fetch              => s_fetch(13,25),
			data_in            => s_data_in(13,25),
			data_out           => s_data_out(13,25),
			out1               => s_out1(13,25),
			out2               => s_out2(13,25),
			lock_lower_row_out => s_locks_lower_out(13,25),
			lock_lower_row_in  => s_locks_lower_in(13,25),
			in1                => s_in1(13,25),
			in2                => s_in2(13,25),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(25)
		);
	s_in1(13,25)            <= s_out1(14,25);
	s_in2(13,25)            <= s_out2(14,26);
	s_locks_lower_in(13,25) <= s_locks_lower_out(14,25);

		normal_cell_13_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,26),
			fetch              => s_fetch(13,26),
			data_in            => s_data_in(13,26),
			data_out           => s_data_out(13,26),
			out1               => s_out1(13,26),
			out2               => s_out2(13,26),
			lock_lower_row_out => s_locks_lower_out(13,26),
			lock_lower_row_in  => s_locks_lower_in(13,26),
			in1                => s_in1(13,26),
			in2                => s_in2(13,26),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(26)
		);
	s_in1(13,26)            <= s_out1(14,26);
	s_in2(13,26)            <= s_out2(14,27);
	s_locks_lower_in(13,26) <= s_locks_lower_out(14,26);

		normal_cell_13_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,27),
			fetch              => s_fetch(13,27),
			data_in            => s_data_in(13,27),
			data_out           => s_data_out(13,27),
			out1               => s_out1(13,27),
			out2               => s_out2(13,27),
			lock_lower_row_out => s_locks_lower_out(13,27),
			lock_lower_row_in  => s_locks_lower_in(13,27),
			in1                => s_in1(13,27),
			in2                => s_in2(13,27),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(27)
		);
	s_in1(13,27)            <= s_out1(14,27);
	s_in2(13,27)            <= s_out2(14,28);
	s_locks_lower_in(13,27) <= s_locks_lower_out(14,27);

		normal_cell_13_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,28),
			fetch              => s_fetch(13,28),
			data_in            => s_data_in(13,28),
			data_out           => s_data_out(13,28),
			out1               => s_out1(13,28),
			out2               => s_out2(13,28),
			lock_lower_row_out => s_locks_lower_out(13,28),
			lock_lower_row_in  => s_locks_lower_in(13,28),
			in1                => s_in1(13,28),
			in2                => s_in2(13,28),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(28)
		);
	s_in1(13,28)            <= s_out1(14,28);
	s_in2(13,28)            <= s_out2(14,29);
	s_locks_lower_in(13,28) <= s_locks_lower_out(14,28);

		normal_cell_13_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,29),
			fetch              => s_fetch(13,29),
			data_in            => s_data_in(13,29),
			data_out           => s_data_out(13,29),
			out1               => s_out1(13,29),
			out2               => s_out2(13,29),
			lock_lower_row_out => s_locks_lower_out(13,29),
			lock_lower_row_in  => s_locks_lower_in(13,29),
			in1                => s_in1(13,29),
			in2                => s_in2(13,29),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(29)
		);
	s_in1(13,29)            <= s_out1(14,29);
	s_in2(13,29)            <= s_out2(14,30);
	s_locks_lower_in(13,29) <= s_locks_lower_out(14,29);

		normal_cell_13_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,30),
			fetch              => s_fetch(13,30),
			data_in            => s_data_in(13,30),
			data_out           => s_data_out(13,30),
			out1               => s_out1(13,30),
			out2               => s_out2(13,30),
			lock_lower_row_out => s_locks_lower_out(13,30),
			lock_lower_row_in  => s_locks_lower_in(13,30),
			in1                => s_in1(13,30),
			in2                => s_in2(13,30),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(30)
		);
	s_in1(13,30)            <= s_out1(14,30);
	s_in2(13,30)            <= s_out2(14,31);
	s_locks_lower_in(13,30) <= s_locks_lower_out(14,30);

		normal_cell_13_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,31),
			fetch              => s_fetch(13,31),
			data_in            => s_data_in(13,31),
			data_out           => s_data_out(13,31),
			out1               => s_out1(13,31),
			out2               => s_out2(13,31),
			lock_lower_row_out => s_locks_lower_out(13,31),
			lock_lower_row_in  => s_locks_lower_in(13,31),
			in1                => s_in1(13,31),
			in2                => s_in2(13,31),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(31)
		);
	s_in1(13,31)            <= s_out1(14,31);
	s_in2(13,31)            <= s_out2(14,32);
	s_locks_lower_in(13,31) <= s_locks_lower_out(14,31);

		normal_cell_13_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,32),
			fetch              => s_fetch(13,32),
			data_in            => s_data_in(13,32),
			data_out           => s_data_out(13,32),
			out1               => s_out1(13,32),
			out2               => s_out2(13,32),
			lock_lower_row_out => s_locks_lower_out(13,32),
			lock_lower_row_in  => s_locks_lower_in(13,32),
			in1                => s_in1(13,32),
			in2                => s_in2(13,32),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(32)
		);
	s_in1(13,32)            <= s_out1(14,32);
	s_in2(13,32)            <= s_out2(14,33);
	s_locks_lower_in(13,32) <= s_locks_lower_out(14,32);

		normal_cell_13_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,33),
			fetch              => s_fetch(13,33),
			data_in            => s_data_in(13,33),
			data_out           => s_data_out(13,33),
			out1               => s_out1(13,33),
			out2               => s_out2(13,33),
			lock_lower_row_out => s_locks_lower_out(13,33),
			lock_lower_row_in  => s_locks_lower_in(13,33),
			in1                => s_in1(13,33),
			in2                => s_in2(13,33),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(33)
		);
	s_in1(13,33)            <= s_out1(14,33);
	s_in2(13,33)            <= s_out2(14,34);
	s_locks_lower_in(13,33) <= s_locks_lower_out(14,33);

		normal_cell_13_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,34),
			fetch              => s_fetch(13,34),
			data_in            => s_data_in(13,34),
			data_out           => s_data_out(13,34),
			out1               => s_out1(13,34),
			out2               => s_out2(13,34),
			lock_lower_row_out => s_locks_lower_out(13,34),
			lock_lower_row_in  => s_locks_lower_in(13,34),
			in1                => s_in1(13,34),
			in2                => s_in2(13,34),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(34)
		);
	s_in1(13,34)            <= s_out1(14,34);
	s_in2(13,34)            <= s_out2(14,35);
	s_locks_lower_in(13,34) <= s_locks_lower_out(14,34);

		normal_cell_13_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,35),
			fetch              => s_fetch(13,35),
			data_in            => s_data_in(13,35),
			data_out           => s_data_out(13,35),
			out1               => s_out1(13,35),
			out2               => s_out2(13,35),
			lock_lower_row_out => s_locks_lower_out(13,35),
			lock_lower_row_in  => s_locks_lower_in(13,35),
			in1                => s_in1(13,35),
			in2                => s_in2(13,35),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(35)
		);
	s_in1(13,35)            <= s_out1(14,35);
	s_in2(13,35)            <= s_out2(14,36);
	s_locks_lower_in(13,35) <= s_locks_lower_out(14,35);

		normal_cell_13_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,36),
			fetch              => s_fetch(13,36),
			data_in            => s_data_in(13,36),
			data_out           => s_data_out(13,36),
			out1               => s_out1(13,36),
			out2               => s_out2(13,36),
			lock_lower_row_out => s_locks_lower_out(13,36),
			lock_lower_row_in  => s_locks_lower_in(13,36),
			in1                => s_in1(13,36),
			in2                => s_in2(13,36),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(36)
		);
	s_in1(13,36)            <= s_out1(14,36);
	s_in2(13,36)            <= s_out2(14,37);
	s_locks_lower_in(13,36) <= s_locks_lower_out(14,36);

		normal_cell_13_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,37),
			fetch              => s_fetch(13,37),
			data_in            => s_data_in(13,37),
			data_out           => s_data_out(13,37),
			out1               => s_out1(13,37),
			out2               => s_out2(13,37),
			lock_lower_row_out => s_locks_lower_out(13,37),
			lock_lower_row_in  => s_locks_lower_in(13,37),
			in1                => s_in1(13,37),
			in2                => s_in2(13,37),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(37)
		);
	s_in1(13,37)            <= s_out1(14,37);
	s_in2(13,37)            <= s_out2(14,38);
	s_locks_lower_in(13,37) <= s_locks_lower_out(14,37);

		normal_cell_13_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,38),
			fetch              => s_fetch(13,38),
			data_in            => s_data_in(13,38),
			data_out           => s_data_out(13,38),
			out1               => s_out1(13,38),
			out2               => s_out2(13,38),
			lock_lower_row_out => s_locks_lower_out(13,38),
			lock_lower_row_in  => s_locks_lower_in(13,38),
			in1                => s_in1(13,38),
			in2                => s_in2(13,38),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(38)
		);
	s_in1(13,38)            <= s_out1(14,38);
	s_in2(13,38)            <= s_out2(14,39);
	s_locks_lower_in(13,38) <= s_locks_lower_out(14,38);

		normal_cell_13_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,39),
			fetch              => s_fetch(13,39),
			data_in            => s_data_in(13,39),
			data_out           => s_data_out(13,39),
			out1               => s_out1(13,39),
			out2               => s_out2(13,39),
			lock_lower_row_out => s_locks_lower_out(13,39),
			lock_lower_row_in  => s_locks_lower_in(13,39),
			in1                => s_in1(13,39),
			in2                => s_in2(13,39),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(39)
		);
	s_in1(13,39)            <= s_out1(14,39);
	s_in2(13,39)            <= s_out2(14,40);
	s_locks_lower_in(13,39) <= s_locks_lower_out(14,39);

		normal_cell_13_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,40),
			fetch              => s_fetch(13,40),
			data_in            => s_data_in(13,40),
			data_out           => s_data_out(13,40),
			out1               => s_out1(13,40),
			out2               => s_out2(13,40),
			lock_lower_row_out => s_locks_lower_out(13,40),
			lock_lower_row_in  => s_locks_lower_in(13,40),
			in1                => s_in1(13,40),
			in2                => s_in2(13,40),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(40)
		);
	s_in1(13,40)            <= s_out1(14,40);
	s_in2(13,40)            <= s_out2(14,41);
	s_locks_lower_in(13,40) <= s_locks_lower_out(14,40);

		normal_cell_13_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,41),
			fetch              => s_fetch(13,41),
			data_in            => s_data_in(13,41),
			data_out           => s_data_out(13,41),
			out1               => s_out1(13,41),
			out2               => s_out2(13,41),
			lock_lower_row_out => s_locks_lower_out(13,41),
			lock_lower_row_in  => s_locks_lower_in(13,41),
			in1                => s_in1(13,41),
			in2                => s_in2(13,41),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(41)
		);
	s_in1(13,41)            <= s_out1(14,41);
	s_in2(13,41)            <= s_out2(14,42);
	s_locks_lower_in(13,41) <= s_locks_lower_out(14,41);

		normal_cell_13_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,42),
			fetch              => s_fetch(13,42),
			data_in            => s_data_in(13,42),
			data_out           => s_data_out(13,42),
			out1               => s_out1(13,42),
			out2               => s_out2(13,42),
			lock_lower_row_out => s_locks_lower_out(13,42),
			lock_lower_row_in  => s_locks_lower_in(13,42),
			in1                => s_in1(13,42),
			in2                => s_in2(13,42),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(42)
		);
	s_in1(13,42)            <= s_out1(14,42);
	s_in2(13,42)            <= s_out2(14,43);
	s_locks_lower_in(13,42) <= s_locks_lower_out(14,42);

		normal_cell_13_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,43),
			fetch              => s_fetch(13,43),
			data_in            => s_data_in(13,43),
			data_out           => s_data_out(13,43),
			out1               => s_out1(13,43),
			out2               => s_out2(13,43),
			lock_lower_row_out => s_locks_lower_out(13,43),
			lock_lower_row_in  => s_locks_lower_in(13,43),
			in1                => s_in1(13,43),
			in2                => s_in2(13,43),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(43)
		);
	s_in1(13,43)            <= s_out1(14,43);
	s_in2(13,43)            <= s_out2(14,44);
	s_locks_lower_in(13,43) <= s_locks_lower_out(14,43);

		normal_cell_13_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,44),
			fetch              => s_fetch(13,44),
			data_in            => s_data_in(13,44),
			data_out           => s_data_out(13,44),
			out1               => s_out1(13,44),
			out2               => s_out2(13,44),
			lock_lower_row_out => s_locks_lower_out(13,44),
			lock_lower_row_in  => s_locks_lower_in(13,44),
			in1                => s_in1(13,44),
			in2                => s_in2(13,44),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(44)
		);
	s_in1(13,44)            <= s_out1(14,44);
	s_in2(13,44)            <= s_out2(14,45);
	s_locks_lower_in(13,44) <= s_locks_lower_out(14,44);

		normal_cell_13_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,45),
			fetch              => s_fetch(13,45),
			data_in            => s_data_in(13,45),
			data_out           => s_data_out(13,45),
			out1               => s_out1(13,45),
			out2               => s_out2(13,45),
			lock_lower_row_out => s_locks_lower_out(13,45),
			lock_lower_row_in  => s_locks_lower_in(13,45),
			in1                => s_in1(13,45),
			in2                => s_in2(13,45),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(45)
		);
	s_in1(13,45)            <= s_out1(14,45);
	s_in2(13,45)            <= s_out2(14,46);
	s_locks_lower_in(13,45) <= s_locks_lower_out(14,45);

		normal_cell_13_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,46),
			fetch              => s_fetch(13,46),
			data_in            => s_data_in(13,46),
			data_out           => s_data_out(13,46),
			out1               => s_out1(13,46),
			out2               => s_out2(13,46),
			lock_lower_row_out => s_locks_lower_out(13,46),
			lock_lower_row_in  => s_locks_lower_in(13,46),
			in1                => s_in1(13,46),
			in2                => s_in2(13,46),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(46)
		);
	s_in1(13,46)            <= s_out1(14,46);
	s_in2(13,46)            <= s_out2(14,47);
	s_locks_lower_in(13,46) <= s_locks_lower_out(14,46);

		normal_cell_13_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,47),
			fetch              => s_fetch(13,47),
			data_in            => s_data_in(13,47),
			data_out           => s_data_out(13,47),
			out1               => s_out1(13,47),
			out2               => s_out2(13,47),
			lock_lower_row_out => s_locks_lower_out(13,47),
			lock_lower_row_in  => s_locks_lower_in(13,47),
			in1                => s_in1(13,47),
			in2                => s_in2(13,47),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(47)
		);
	s_in1(13,47)            <= s_out1(14,47);
	s_in2(13,47)            <= s_out2(14,48);
	s_locks_lower_in(13,47) <= s_locks_lower_out(14,47);

		normal_cell_13_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,48),
			fetch              => s_fetch(13,48),
			data_in            => s_data_in(13,48),
			data_out           => s_data_out(13,48),
			out1               => s_out1(13,48),
			out2               => s_out2(13,48),
			lock_lower_row_out => s_locks_lower_out(13,48),
			lock_lower_row_in  => s_locks_lower_in(13,48),
			in1                => s_in1(13,48),
			in2                => s_in2(13,48),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(48)
		);
	s_in1(13,48)            <= s_out1(14,48);
	s_in2(13,48)            <= s_out2(14,49);
	s_locks_lower_in(13,48) <= s_locks_lower_out(14,48);

		normal_cell_13_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,49),
			fetch              => s_fetch(13,49),
			data_in            => s_data_in(13,49),
			data_out           => s_data_out(13,49),
			out1               => s_out1(13,49),
			out2               => s_out2(13,49),
			lock_lower_row_out => s_locks_lower_out(13,49),
			lock_lower_row_in  => s_locks_lower_in(13,49),
			in1                => s_in1(13,49),
			in2                => s_in2(13,49),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(49)
		);
	s_in1(13,49)            <= s_out1(14,49);
	s_in2(13,49)            <= s_out2(14,50);
	s_locks_lower_in(13,49) <= s_locks_lower_out(14,49);

		normal_cell_13_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,50),
			fetch              => s_fetch(13,50),
			data_in            => s_data_in(13,50),
			data_out           => s_data_out(13,50),
			out1               => s_out1(13,50),
			out2               => s_out2(13,50),
			lock_lower_row_out => s_locks_lower_out(13,50),
			lock_lower_row_in  => s_locks_lower_in(13,50),
			in1                => s_in1(13,50),
			in2                => s_in2(13,50),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(50)
		);
	s_in1(13,50)            <= s_out1(14,50);
	s_in2(13,50)            <= s_out2(14,51);
	s_locks_lower_in(13,50) <= s_locks_lower_out(14,50);

		normal_cell_13_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,51),
			fetch              => s_fetch(13,51),
			data_in            => s_data_in(13,51),
			data_out           => s_data_out(13,51),
			out1               => s_out1(13,51),
			out2               => s_out2(13,51),
			lock_lower_row_out => s_locks_lower_out(13,51),
			lock_lower_row_in  => s_locks_lower_in(13,51),
			in1                => s_in1(13,51),
			in2                => s_in2(13,51),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(51)
		);
	s_in1(13,51)            <= s_out1(14,51);
	s_in2(13,51)            <= s_out2(14,52);
	s_locks_lower_in(13,51) <= s_locks_lower_out(14,51);

		normal_cell_13_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,52),
			fetch              => s_fetch(13,52),
			data_in            => s_data_in(13,52),
			data_out           => s_data_out(13,52),
			out1               => s_out1(13,52),
			out2               => s_out2(13,52),
			lock_lower_row_out => s_locks_lower_out(13,52),
			lock_lower_row_in  => s_locks_lower_in(13,52),
			in1                => s_in1(13,52),
			in2                => s_in2(13,52),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(52)
		);
	s_in1(13,52)            <= s_out1(14,52);
	s_in2(13,52)            <= s_out2(14,53);
	s_locks_lower_in(13,52) <= s_locks_lower_out(14,52);

		normal_cell_13_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,53),
			fetch              => s_fetch(13,53),
			data_in            => s_data_in(13,53),
			data_out           => s_data_out(13,53),
			out1               => s_out1(13,53),
			out2               => s_out2(13,53),
			lock_lower_row_out => s_locks_lower_out(13,53),
			lock_lower_row_in  => s_locks_lower_in(13,53),
			in1                => s_in1(13,53),
			in2                => s_in2(13,53),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(53)
		);
	s_in1(13,53)            <= s_out1(14,53);
	s_in2(13,53)            <= s_out2(14,54);
	s_locks_lower_in(13,53) <= s_locks_lower_out(14,53);

		normal_cell_13_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,54),
			fetch              => s_fetch(13,54),
			data_in            => s_data_in(13,54),
			data_out           => s_data_out(13,54),
			out1               => s_out1(13,54),
			out2               => s_out2(13,54),
			lock_lower_row_out => s_locks_lower_out(13,54),
			lock_lower_row_in  => s_locks_lower_in(13,54),
			in1                => s_in1(13,54),
			in2                => s_in2(13,54),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(54)
		);
	s_in1(13,54)            <= s_out1(14,54);
	s_in2(13,54)            <= s_out2(14,55);
	s_locks_lower_in(13,54) <= s_locks_lower_out(14,54);

		normal_cell_13_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,55),
			fetch              => s_fetch(13,55),
			data_in            => s_data_in(13,55),
			data_out           => s_data_out(13,55),
			out1               => s_out1(13,55),
			out2               => s_out2(13,55),
			lock_lower_row_out => s_locks_lower_out(13,55),
			lock_lower_row_in  => s_locks_lower_in(13,55),
			in1                => s_in1(13,55),
			in2                => s_in2(13,55),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(55)
		);
	s_in1(13,55)            <= s_out1(14,55);
	s_in2(13,55)            <= s_out2(14,56);
	s_locks_lower_in(13,55) <= s_locks_lower_out(14,55);

		normal_cell_13_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,56),
			fetch              => s_fetch(13,56),
			data_in            => s_data_in(13,56),
			data_out           => s_data_out(13,56),
			out1               => s_out1(13,56),
			out2               => s_out2(13,56),
			lock_lower_row_out => s_locks_lower_out(13,56),
			lock_lower_row_in  => s_locks_lower_in(13,56),
			in1                => s_in1(13,56),
			in2                => s_in2(13,56),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(56)
		);
	s_in1(13,56)            <= s_out1(14,56);
	s_in2(13,56)            <= s_out2(14,57);
	s_locks_lower_in(13,56) <= s_locks_lower_out(14,56);

		normal_cell_13_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,57),
			fetch              => s_fetch(13,57),
			data_in            => s_data_in(13,57),
			data_out           => s_data_out(13,57),
			out1               => s_out1(13,57),
			out2               => s_out2(13,57),
			lock_lower_row_out => s_locks_lower_out(13,57),
			lock_lower_row_in  => s_locks_lower_in(13,57),
			in1                => s_in1(13,57),
			in2                => s_in2(13,57),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(57)
		);
	s_in1(13,57)            <= s_out1(14,57);
	s_in2(13,57)            <= s_out2(14,58);
	s_locks_lower_in(13,57) <= s_locks_lower_out(14,57);

		normal_cell_13_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,58),
			fetch              => s_fetch(13,58),
			data_in            => s_data_in(13,58),
			data_out           => s_data_out(13,58),
			out1               => s_out1(13,58),
			out2               => s_out2(13,58),
			lock_lower_row_out => s_locks_lower_out(13,58),
			lock_lower_row_in  => s_locks_lower_in(13,58),
			in1                => s_in1(13,58),
			in2                => s_in2(13,58),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(58)
		);
	s_in1(13,58)            <= s_out1(14,58);
	s_in2(13,58)            <= s_out2(14,59);
	s_locks_lower_in(13,58) <= s_locks_lower_out(14,58);

		normal_cell_13_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,59),
			fetch              => s_fetch(13,59),
			data_in            => s_data_in(13,59),
			data_out           => s_data_out(13,59),
			out1               => s_out1(13,59),
			out2               => s_out2(13,59),
			lock_lower_row_out => s_locks_lower_out(13,59),
			lock_lower_row_in  => s_locks_lower_in(13,59),
			in1                => s_in1(13,59),
			in2                => s_in2(13,59),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(59)
		);
	s_in1(13,59)            <= s_out1(14,59);
	s_in2(13,59)            <= s_out2(14,60);
	s_locks_lower_in(13,59) <= s_locks_lower_out(14,59);

		last_col_cell_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(13,60),
			fetch              => s_fetch(13,60),
			data_in            => s_data_in(13,60),
			data_out           => s_data_out(13,60),
			out1               => s_out1(13,60),
			out2               => s_out2(13,60),
			lock_lower_row_out => s_locks_lower_out(13,60),
			lock_lower_row_in  => s_locks_lower_in(13,60),
			in1                => s_in1(13,60),
			in2                => (others => '0'),
			lock_row           => s_locks(13),
			piv_found          => s_piv_found,
			row_data           => s_row_data(13),
			col_data           => s_col_data(60)
		);
	s_in1(13,60)            <= s_out1(14,60);
	s_locks_lower_in(13,60) <= s_locks_lower_out(14,60);

		normal_cell_14_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,1),
			fetch              => s_fetch(14,1),
			data_in            => s_data_in(14,1),
			data_out           => s_data_out(14,1),
			out1               => s_out1(14,1),
			out2               => s_out2(14,1),
			lock_lower_row_out => s_locks_lower_out(14,1),
			lock_lower_row_in  => s_locks_lower_in(14,1),
			in1                => s_in1(14,1),
			in2                => s_in2(14,1),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(1)
		);
	s_in1(14,1)            <= s_out1(15,1);
	s_in2(14,1)            <= s_out2(15,2);
	s_locks_lower_in(14,1) <= s_locks_lower_out(15,1);

		normal_cell_14_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,2),
			fetch              => s_fetch(14,2),
			data_in            => s_data_in(14,2),
			data_out           => s_data_out(14,2),
			out1               => s_out1(14,2),
			out2               => s_out2(14,2),
			lock_lower_row_out => s_locks_lower_out(14,2),
			lock_lower_row_in  => s_locks_lower_in(14,2),
			in1                => s_in1(14,2),
			in2                => s_in2(14,2),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(2)
		);
	s_in1(14,2)            <= s_out1(15,2);
	s_in2(14,2)            <= s_out2(15,3);
	s_locks_lower_in(14,2) <= s_locks_lower_out(15,2);

		normal_cell_14_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,3),
			fetch              => s_fetch(14,3),
			data_in            => s_data_in(14,3),
			data_out           => s_data_out(14,3),
			out1               => s_out1(14,3),
			out2               => s_out2(14,3),
			lock_lower_row_out => s_locks_lower_out(14,3),
			lock_lower_row_in  => s_locks_lower_in(14,3),
			in1                => s_in1(14,3),
			in2                => s_in2(14,3),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(3)
		);
	s_in1(14,3)            <= s_out1(15,3);
	s_in2(14,3)            <= s_out2(15,4);
	s_locks_lower_in(14,3) <= s_locks_lower_out(15,3);

		normal_cell_14_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,4),
			fetch              => s_fetch(14,4),
			data_in            => s_data_in(14,4),
			data_out           => s_data_out(14,4),
			out1               => s_out1(14,4),
			out2               => s_out2(14,4),
			lock_lower_row_out => s_locks_lower_out(14,4),
			lock_lower_row_in  => s_locks_lower_in(14,4),
			in1                => s_in1(14,4),
			in2                => s_in2(14,4),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(4)
		);
	s_in1(14,4)            <= s_out1(15,4);
	s_in2(14,4)            <= s_out2(15,5);
	s_locks_lower_in(14,4) <= s_locks_lower_out(15,4);

		normal_cell_14_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,5),
			fetch              => s_fetch(14,5),
			data_in            => s_data_in(14,5),
			data_out           => s_data_out(14,5),
			out1               => s_out1(14,5),
			out2               => s_out2(14,5),
			lock_lower_row_out => s_locks_lower_out(14,5),
			lock_lower_row_in  => s_locks_lower_in(14,5),
			in1                => s_in1(14,5),
			in2                => s_in2(14,5),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(5)
		);
	s_in1(14,5)            <= s_out1(15,5);
	s_in2(14,5)            <= s_out2(15,6);
	s_locks_lower_in(14,5) <= s_locks_lower_out(15,5);

		normal_cell_14_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,6),
			fetch              => s_fetch(14,6),
			data_in            => s_data_in(14,6),
			data_out           => s_data_out(14,6),
			out1               => s_out1(14,6),
			out2               => s_out2(14,6),
			lock_lower_row_out => s_locks_lower_out(14,6),
			lock_lower_row_in  => s_locks_lower_in(14,6),
			in1                => s_in1(14,6),
			in2                => s_in2(14,6),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(6)
		);
	s_in1(14,6)            <= s_out1(15,6);
	s_in2(14,6)            <= s_out2(15,7);
	s_locks_lower_in(14,6) <= s_locks_lower_out(15,6);

		normal_cell_14_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,7),
			fetch              => s_fetch(14,7),
			data_in            => s_data_in(14,7),
			data_out           => s_data_out(14,7),
			out1               => s_out1(14,7),
			out2               => s_out2(14,7),
			lock_lower_row_out => s_locks_lower_out(14,7),
			lock_lower_row_in  => s_locks_lower_in(14,7),
			in1                => s_in1(14,7),
			in2                => s_in2(14,7),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(7)
		);
	s_in1(14,7)            <= s_out1(15,7);
	s_in2(14,7)            <= s_out2(15,8);
	s_locks_lower_in(14,7) <= s_locks_lower_out(15,7);

		normal_cell_14_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,8),
			fetch              => s_fetch(14,8),
			data_in            => s_data_in(14,8),
			data_out           => s_data_out(14,8),
			out1               => s_out1(14,8),
			out2               => s_out2(14,8),
			lock_lower_row_out => s_locks_lower_out(14,8),
			lock_lower_row_in  => s_locks_lower_in(14,8),
			in1                => s_in1(14,8),
			in2                => s_in2(14,8),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(8)
		);
	s_in1(14,8)            <= s_out1(15,8);
	s_in2(14,8)            <= s_out2(15,9);
	s_locks_lower_in(14,8) <= s_locks_lower_out(15,8);

		normal_cell_14_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,9),
			fetch              => s_fetch(14,9),
			data_in            => s_data_in(14,9),
			data_out           => s_data_out(14,9),
			out1               => s_out1(14,9),
			out2               => s_out2(14,9),
			lock_lower_row_out => s_locks_lower_out(14,9),
			lock_lower_row_in  => s_locks_lower_in(14,9),
			in1                => s_in1(14,9),
			in2                => s_in2(14,9),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(9)
		);
	s_in1(14,9)            <= s_out1(15,9);
	s_in2(14,9)            <= s_out2(15,10);
	s_locks_lower_in(14,9) <= s_locks_lower_out(15,9);

		normal_cell_14_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,10),
			fetch              => s_fetch(14,10),
			data_in            => s_data_in(14,10),
			data_out           => s_data_out(14,10),
			out1               => s_out1(14,10),
			out2               => s_out2(14,10),
			lock_lower_row_out => s_locks_lower_out(14,10),
			lock_lower_row_in  => s_locks_lower_in(14,10),
			in1                => s_in1(14,10),
			in2                => s_in2(14,10),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(10)
		);
	s_in1(14,10)            <= s_out1(15,10);
	s_in2(14,10)            <= s_out2(15,11);
	s_locks_lower_in(14,10) <= s_locks_lower_out(15,10);

		normal_cell_14_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,11),
			fetch              => s_fetch(14,11),
			data_in            => s_data_in(14,11),
			data_out           => s_data_out(14,11),
			out1               => s_out1(14,11),
			out2               => s_out2(14,11),
			lock_lower_row_out => s_locks_lower_out(14,11),
			lock_lower_row_in  => s_locks_lower_in(14,11),
			in1                => s_in1(14,11),
			in2                => s_in2(14,11),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(11)
		);
	s_in1(14,11)            <= s_out1(15,11);
	s_in2(14,11)            <= s_out2(15,12);
	s_locks_lower_in(14,11) <= s_locks_lower_out(15,11);

		normal_cell_14_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,12),
			fetch              => s_fetch(14,12),
			data_in            => s_data_in(14,12),
			data_out           => s_data_out(14,12),
			out1               => s_out1(14,12),
			out2               => s_out2(14,12),
			lock_lower_row_out => s_locks_lower_out(14,12),
			lock_lower_row_in  => s_locks_lower_in(14,12),
			in1                => s_in1(14,12),
			in2                => s_in2(14,12),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(12)
		);
	s_in1(14,12)            <= s_out1(15,12);
	s_in2(14,12)            <= s_out2(15,13);
	s_locks_lower_in(14,12) <= s_locks_lower_out(15,12);

		normal_cell_14_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,13),
			fetch              => s_fetch(14,13),
			data_in            => s_data_in(14,13),
			data_out           => s_data_out(14,13),
			out1               => s_out1(14,13),
			out2               => s_out2(14,13),
			lock_lower_row_out => s_locks_lower_out(14,13),
			lock_lower_row_in  => s_locks_lower_in(14,13),
			in1                => s_in1(14,13),
			in2                => s_in2(14,13),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(13)
		);
	s_in1(14,13)            <= s_out1(15,13);
	s_in2(14,13)            <= s_out2(15,14);
	s_locks_lower_in(14,13) <= s_locks_lower_out(15,13);

		normal_cell_14_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,14),
			fetch              => s_fetch(14,14),
			data_in            => s_data_in(14,14),
			data_out           => s_data_out(14,14),
			out1               => s_out1(14,14),
			out2               => s_out2(14,14),
			lock_lower_row_out => s_locks_lower_out(14,14),
			lock_lower_row_in  => s_locks_lower_in(14,14),
			in1                => s_in1(14,14),
			in2                => s_in2(14,14),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(14)
		);
	s_in1(14,14)            <= s_out1(15,14);
	s_in2(14,14)            <= s_out2(15,15);
	s_locks_lower_in(14,14) <= s_locks_lower_out(15,14);

		normal_cell_14_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,15),
			fetch              => s_fetch(14,15),
			data_in            => s_data_in(14,15),
			data_out           => s_data_out(14,15),
			out1               => s_out1(14,15),
			out2               => s_out2(14,15),
			lock_lower_row_out => s_locks_lower_out(14,15),
			lock_lower_row_in  => s_locks_lower_in(14,15),
			in1                => s_in1(14,15),
			in2                => s_in2(14,15),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(15)
		);
	s_in1(14,15)            <= s_out1(15,15);
	s_in2(14,15)            <= s_out2(15,16);
	s_locks_lower_in(14,15) <= s_locks_lower_out(15,15);

		normal_cell_14_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,16),
			fetch              => s_fetch(14,16),
			data_in            => s_data_in(14,16),
			data_out           => s_data_out(14,16),
			out1               => s_out1(14,16),
			out2               => s_out2(14,16),
			lock_lower_row_out => s_locks_lower_out(14,16),
			lock_lower_row_in  => s_locks_lower_in(14,16),
			in1                => s_in1(14,16),
			in2                => s_in2(14,16),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(16)
		);
	s_in1(14,16)            <= s_out1(15,16);
	s_in2(14,16)            <= s_out2(15,17);
	s_locks_lower_in(14,16) <= s_locks_lower_out(15,16);

		normal_cell_14_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,17),
			fetch              => s_fetch(14,17),
			data_in            => s_data_in(14,17),
			data_out           => s_data_out(14,17),
			out1               => s_out1(14,17),
			out2               => s_out2(14,17),
			lock_lower_row_out => s_locks_lower_out(14,17),
			lock_lower_row_in  => s_locks_lower_in(14,17),
			in1                => s_in1(14,17),
			in2                => s_in2(14,17),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(17)
		);
	s_in1(14,17)            <= s_out1(15,17);
	s_in2(14,17)            <= s_out2(15,18);
	s_locks_lower_in(14,17) <= s_locks_lower_out(15,17);

		normal_cell_14_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,18),
			fetch              => s_fetch(14,18),
			data_in            => s_data_in(14,18),
			data_out           => s_data_out(14,18),
			out1               => s_out1(14,18),
			out2               => s_out2(14,18),
			lock_lower_row_out => s_locks_lower_out(14,18),
			lock_lower_row_in  => s_locks_lower_in(14,18),
			in1                => s_in1(14,18),
			in2                => s_in2(14,18),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(18)
		);
	s_in1(14,18)            <= s_out1(15,18);
	s_in2(14,18)            <= s_out2(15,19);
	s_locks_lower_in(14,18) <= s_locks_lower_out(15,18);

		normal_cell_14_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,19),
			fetch              => s_fetch(14,19),
			data_in            => s_data_in(14,19),
			data_out           => s_data_out(14,19),
			out1               => s_out1(14,19),
			out2               => s_out2(14,19),
			lock_lower_row_out => s_locks_lower_out(14,19),
			lock_lower_row_in  => s_locks_lower_in(14,19),
			in1                => s_in1(14,19),
			in2                => s_in2(14,19),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(19)
		);
	s_in1(14,19)            <= s_out1(15,19);
	s_in2(14,19)            <= s_out2(15,20);
	s_locks_lower_in(14,19) <= s_locks_lower_out(15,19);

		normal_cell_14_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,20),
			fetch              => s_fetch(14,20),
			data_in            => s_data_in(14,20),
			data_out           => s_data_out(14,20),
			out1               => s_out1(14,20),
			out2               => s_out2(14,20),
			lock_lower_row_out => s_locks_lower_out(14,20),
			lock_lower_row_in  => s_locks_lower_in(14,20),
			in1                => s_in1(14,20),
			in2                => s_in2(14,20),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(20)
		);
	s_in1(14,20)            <= s_out1(15,20);
	s_in2(14,20)            <= s_out2(15,21);
	s_locks_lower_in(14,20) <= s_locks_lower_out(15,20);

		normal_cell_14_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,21),
			fetch              => s_fetch(14,21),
			data_in            => s_data_in(14,21),
			data_out           => s_data_out(14,21),
			out1               => s_out1(14,21),
			out2               => s_out2(14,21),
			lock_lower_row_out => s_locks_lower_out(14,21),
			lock_lower_row_in  => s_locks_lower_in(14,21),
			in1                => s_in1(14,21),
			in2                => s_in2(14,21),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(21)
		);
	s_in1(14,21)            <= s_out1(15,21);
	s_in2(14,21)            <= s_out2(15,22);
	s_locks_lower_in(14,21) <= s_locks_lower_out(15,21);

		normal_cell_14_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,22),
			fetch              => s_fetch(14,22),
			data_in            => s_data_in(14,22),
			data_out           => s_data_out(14,22),
			out1               => s_out1(14,22),
			out2               => s_out2(14,22),
			lock_lower_row_out => s_locks_lower_out(14,22),
			lock_lower_row_in  => s_locks_lower_in(14,22),
			in1                => s_in1(14,22),
			in2                => s_in2(14,22),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(22)
		);
	s_in1(14,22)            <= s_out1(15,22);
	s_in2(14,22)            <= s_out2(15,23);
	s_locks_lower_in(14,22) <= s_locks_lower_out(15,22);

		normal_cell_14_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,23),
			fetch              => s_fetch(14,23),
			data_in            => s_data_in(14,23),
			data_out           => s_data_out(14,23),
			out1               => s_out1(14,23),
			out2               => s_out2(14,23),
			lock_lower_row_out => s_locks_lower_out(14,23),
			lock_lower_row_in  => s_locks_lower_in(14,23),
			in1                => s_in1(14,23),
			in2                => s_in2(14,23),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(23)
		);
	s_in1(14,23)            <= s_out1(15,23);
	s_in2(14,23)            <= s_out2(15,24);
	s_locks_lower_in(14,23) <= s_locks_lower_out(15,23);

		normal_cell_14_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,24),
			fetch              => s_fetch(14,24),
			data_in            => s_data_in(14,24),
			data_out           => s_data_out(14,24),
			out1               => s_out1(14,24),
			out2               => s_out2(14,24),
			lock_lower_row_out => s_locks_lower_out(14,24),
			lock_lower_row_in  => s_locks_lower_in(14,24),
			in1                => s_in1(14,24),
			in2                => s_in2(14,24),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(24)
		);
	s_in1(14,24)            <= s_out1(15,24);
	s_in2(14,24)            <= s_out2(15,25);
	s_locks_lower_in(14,24) <= s_locks_lower_out(15,24);

		normal_cell_14_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,25),
			fetch              => s_fetch(14,25),
			data_in            => s_data_in(14,25),
			data_out           => s_data_out(14,25),
			out1               => s_out1(14,25),
			out2               => s_out2(14,25),
			lock_lower_row_out => s_locks_lower_out(14,25),
			lock_lower_row_in  => s_locks_lower_in(14,25),
			in1                => s_in1(14,25),
			in2                => s_in2(14,25),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(25)
		);
	s_in1(14,25)            <= s_out1(15,25);
	s_in2(14,25)            <= s_out2(15,26);
	s_locks_lower_in(14,25) <= s_locks_lower_out(15,25);

		normal_cell_14_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,26),
			fetch              => s_fetch(14,26),
			data_in            => s_data_in(14,26),
			data_out           => s_data_out(14,26),
			out1               => s_out1(14,26),
			out2               => s_out2(14,26),
			lock_lower_row_out => s_locks_lower_out(14,26),
			lock_lower_row_in  => s_locks_lower_in(14,26),
			in1                => s_in1(14,26),
			in2                => s_in2(14,26),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(26)
		);
	s_in1(14,26)            <= s_out1(15,26);
	s_in2(14,26)            <= s_out2(15,27);
	s_locks_lower_in(14,26) <= s_locks_lower_out(15,26);

		normal_cell_14_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,27),
			fetch              => s_fetch(14,27),
			data_in            => s_data_in(14,27),
			data_out           => s_data_out(14,27),
			out1               => s_out1(14,27),
			out2               => s_out2(14,27),
			lock_lower_row_out => s_locks_lower_out(14,27),
			lock_lower_row_in  => s_locks_lower_in(14,27),
			in1                => s_in1(14,27),
			in2                => s_in2(14,27),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(27)
		);
	s_in1(14,27)            <= s_out1(15,27);
	s_in2(14,27)            <= s_out2(15,28);
	s_locks_lower_in(14,27) <= s_locks_lower_out(15,27);

		normal_cell_14_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,28),
			fetch              => s_fetch(14,28),
			data_in            => s_data_in(14,28),
			data_out           => s_data_out(14,28),
			out1               => s_out1(14,28),
			out2               => s_out2(14,28),
			lock_lower_row_out => s_locks_lower_out(14,28),
			lock_lower_row_in  => s_locks_lower_in(14,28),
			in1                => s_in1(14,28),
			in2                => s_in2(14,28),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(28)
		);
	s_in1(14,28)            <= s_out1(15,28);
	s_in2(14,28)            <= s_out2(15,29);
	s_locks_lower_in(14,28) <= s_locks_lower_out(15,28);

		normal_cell_14_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,29),
			fetch              => s_fetch(14,29),
			data_in            => s_data_in(14,29),
			data_out           => s_data_out(14,29),
			out1               => s_out1(14,29),
			out2               => s_out2(14,29),
			lock_lower_row_out => s_locks_lower_out(14,29),
			lock_lower_row_in  => s_locks_lower_in(14,29),
			in1                => s_in1(14,29),
			in2                => s_in2(14,29),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(29)
		);
	s_in1(14,29)            <= s_out1(15,29);
	s_in2(14,29)            <= s_out2(15,30);
	s_locks_lower_in(14,29) <= s_locks_lower_out(15,29);

		normal_cell_14_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,30),
			fetch              => s_fetch(14,30),
			data_in            => s_data_in(14,30),
			data_out           => s_data_out(14,30),
			out1               => s_out1(14,30),
			out2               => s_out2(14,30),
			lock_lower_row_out => s_locks_lower_out(14,30),
			lock_lower_row_in  => s_locks_lower_in(14,30),
			in1                => s_in1(14,30),
			in2                => s_in2(14,30),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(30)
		);
	s_in1(14,30)            <= s_out1(15,30);
	s_in2(14,30)            <= s_out2(15,31);
	s_locks_lower_in(14,30) <= s_locks_lower_out(15,30);

		normal_cell_14_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,31),
			fetch              => s_fetch(14,31),
			data_in            => s_data_in(14,31),
			data_out           => s_data_out(14,31),
			out1               => s_out1(14,31),
			out2               => s_out2(14,31),
			lock_lower_row_out => s_locks_lower_out(14,31),
			lock_lower_row_in  => s_locks_lower_in(14,31),
			in1                => s_in1(14,31),
			in2                => s_in2(14,31),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(31)
		);
	s_in1(14,31)            <= s_out1(15,31);
	s_in2(14,31)            <= s_out2(15,32);
	s_locks_lower_in(14,31) <= s_locks_lower_out(15,31);

		normal_cell_14_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,32),
			fetch              => s_fetch(14,32),
			data_in            => s_data_in(14,32),
			data_out           => s_data_out(14,32),
			out1               => s_out1(14,32),
			out2               => s_out2(14,32),
			lock_lower_row_out => s_locks_lower_out(14,32),
			lock_lower_row_in  => s_locks_lower_in(14,32),
			in1                => s_in1(14,32),
			in2                => s_in2(14,32),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(32)
		);
	s_in1(14,32)            <= s_out1(15,32);
	s_in2(14,32)            <= s_out2(15,33);
	s_locks_lower_in(14,32) <= s_locks_lower_out(15,32);

		normal_cell_14_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,33),
			fetch              => s_fetch(14,33),
			data_in            => s_data_in(14,33),
			data_out           => s_data_out(14,33),
			out1               => s_out1(14,33),
			out2               => s_out2(14,33),
			lock_lower_row_out => s_locks_lower_out(14,33),
			lock_lower_row_in  => s_locks_lower_in(14,33),
			in1                => s_in1(14,33),
			in2                => s_in2(14,33),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(33)
		);
	s_in1(14,33)            <= s_out1(15,33);
	s_in2(14,33)            <= s_out2(15,34);
	s_locks_lower_in(14,33) <= s_locks_lower_out(15,33);

		normal_cell_14_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,34),
			fetch              => s_fetch(14,34),
			data_in            => s_data_in(14,34),
			data_out           => s_data_out(14,34),
			out1               => s_out1(14,34),
			out2               => s_out2(14,34),
			lock_lower_row_out => s_locks_lower_out(14,34),
			lock_lower_row_in  => s_locks_lower_in(14,34),
			in1                => s_in1(14,34),
			in2                => s_in2(14,34),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(34)
		);
	s_in1(14,34)            <= s_out1(15,34);
	s_in2(14,34)            <= s_out2(15,35);
	s_locks_lower_in(14,34) <= s_locks_lower_out(15,34);

		normal_cell_14_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,35),
			fetch              => s_fetch(14,35),
			data_in            => s_data_in(14,35),
			data_out           => s_data_out(14,35),
			out1               => s_out1(14,35),
			out2               => s_out2(14,35),
			lock_lower_row_out => s_locks_lower_out(14,35),
			lock_lower_row_in  => s_locks_lower_in(14,35),
			in1                => s_in1(14,35),
			in2                => s_in2(14,35),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(35)
		);
	s_in1(14,35)            <= s_out1(15,35);
	s_in2(14,35)            <= s_out2(15,36);
	s_locks_lower_in(14,35) <= s_locks_lower_out(15,35);

		normal_cell_14_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,36),
			fetch              => s_fetch(14,36),
			data_in            => s_data_in(14,36),
			data_out           => s_data_out(14,36),
			out1               => s_out1(14,36),
			out2               => s_out2(14,36),
			lock_lower_row_out => s_locks_lower_out(14,36),
			lock_lower_row_in  => s_locks_lower_in(14,36),
			in1                => s_in1(14,36),
			in2                => s_in2(14,36),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(36)
		);
	s_in1(14,36)            <= s_out1(15,36);
	s_in2(14,36)            <= s_out2(15,37);
	s_locks_lower_in(14,36) <= s_locks_lower_out(15,36);

		normal_cell_14_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,37),
			fetch              => s_fetch(14,37),
			data_in            => s_data_in(14,37),
			data_out           => s_data_out(14,37),
			out1               => s_out1(14,37),
			out2               => s_out2(14,37),
			lock_lower_row_out => s_locks_lower_out(14,37),
			lock_lower_row_in  => s_locks_lower_in(14,37),
			in1                => s_in1(14,37),
			in2                => s_in2(14,37),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(37)
		);
	s_in1(14,37)            <= s_out1(15,37);
	s_in2(14,37)            <= s_out2(15,38);
	s_locks_lower_in(14,37) <= s_locks_lower_out(15,37);

		normal_cell_14_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,38),
			fetch              => s_fetch(14,38),
			data_in            => s_data_in(14,38),
			data_out           => s_data_out(14,38),
			out1               => s_out1(14,38),
			out2               => s_out2(14,38),
			lock_lower_row_out => s_locks_lower_out(14,38),
			lock_lower_row_in  => s_locks_lower_in(14,38),
			in1                => s_in1(14,38),
			in2                => s_in2(14,38),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(38)
		);
	s_in1(14,38)            <= s_out1(15,38);
	s_in2(14,38)            <= s_out2(15,39);
	s_locks_lower_in(14,38) <= s_locks_lower_out(15,38);

		normal_cell_14_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,39),
			fetch              => s_fetch(14,39),
			data_in            => s_data_in(14,39),
			data_out           => s_data_out(14,39),
			out1               => s_out1(14,39),
			out2               => s_out2(14,39),
			lock_lower_row_out => s_locks_lower_out(14,39),
			lock_lower_row_in  => s_locks_lower_in(14,39),
			in1                => s_in1(14,39),
			in2                => s_in2(14,39),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(39)
		);
	s_in1(14,39)            <= s_out1(15,39);
	s_in2(14,39)            <= s_out2(15,40);
	s_locks_lower_in(14,39) <= s_locks_lower_out(15,39);

		normal_cell_14_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,40),
			fetch              => s_fetch(14,40),
			data_in            => s_data_in(14,40),
			data_out           => s_data_out(14,40),
			out1               => s_out1(14,40),
			out2               => s_out2(14,40),
			lock_lower_row_out => s_locks_lower_out(14,40),
			lock_lower_row_in  => s_locks_lower_in(14,40),
			in1                => s_in1(14,40),
			in2                => s_in2(14,40),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(40)
		);
	s_in1(14,40)            <= s_out1(15,40);
	s_in2(14,40)            <= s_out2(15,41);
	s_locks_lower_in(14,40) <= s_locks_lower_out(15,40);

		normal_cell_14_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,41),
			fetch              => s_fetch(14,41),
			data_in            => s_data_in(14,41),
			data_out           => s_data_out(14,41),
			out1               => s_out1(14,41),
			out2               => s_out2(14,41),
			lock_lower_row_out => s_locks_lower_out(14,41),
			lock_lower_row_in  => s_locks_lower_in(14,41),
			in1                => s_in1(14,41),
			in2                => s_in2(14,41),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(41)
		);
	s_in1(14,41)            <= s_out1(15,41);
	s_in2(14,41)            <= s_out2(15,42);
	s_locks_lower_in(14,41) <= s_locks_lower_out(15,41);

		normal_cell_14_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,42),
			fetch              => s_fetch(14,42),
			data_in            => s_data_in(14,42),
			data_out           => s_data_out(14,42),
			out1               => s_out1(14,42),
			out2               => s_out2(14,42),
			lock_lower_row_out => s_locks_lower_out(14,42),
			lock_lower_row_in  => s_locks_lower_in(14,42),
			in1                => s_in1(14,42),
			in2                => s_in2(14,42),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(42)
		);
	s_in1(14,42)            <= s_out1(15,42);
	s_in2(14,42)            <= s_out2(15,43);
	s_locks_lower_in(14,42) <= s_locks_lower_out(15,42);

		normal_cell_14_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,43),
			fetch              => s_fetch(14,43),
			data_in            => s_data_in(14,43),
			data_out           => s_data_out(14,43),
			out1               => s_out1(14,43),
			out2               => s_out2(14,43),
			lock_lower_row_out => s_locks_lower_out(14,43),
			lock_lower_row_in  => s_locks_lower_in(14,43),
			in1                => s_in1(14,43),
			in2                => s_in2(14,43),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(43)
		);
	s_in1(14,43)            <= s_out1(15,43);
	s_in2(14,43)            <= s_out2(15,44);
	s_locks_lower_in(14,43) <= s_locks_lower_out(15,43);

		normal_cell_14_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,44),
			fetch              => s_fetch(14,44),
			data_in            => s_data_in(14,44),
			data_out           => s_data_out(14,44),
			out1               => s_out1(14,44),
			out2               => s_out2(14,44),
			lock_lower_row_out => s_locks_lower_out(14,44),
			lock_lower_row_in  => s_locks_lower_in(14,44),
			in1                => s_in1(14,44),
			in2                => s_in2(14,44),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(44)
		);
	s_in1(14,44)            <= s_out1(15,44);
	s_in2(14,44)            <= s_out2(15,45);
	s_locks_lower_in(14,44) <= s_locks_lower_out(15,44);

		normal_cell_14_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,45),
			fetch              => s_fetch(14,45),
			data_in            => s_data_in(14,45),
			data_out           => s_data_out(14,45),
			out1               => s_out1(14,45),
			out2               => s_out2(14,45),
			lock_lower_row_out => s_locks_lower_out(14,45),
			lock_lower_row_in  => s_locks_lower_in(14,45),
			in1                => s_in1(14,45),
			in2                => s_in2(14,45),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(45)
		);
	s_in1(14,45)            <= s_out1(15,45);
	s_in2(14,45)            <= s_out2(15,46);
	s_locks_lower_in(14,45) <= s_locks_lower_out(15,45);

		normal_cell_14_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,46),
			fetch              => s_fetch(14,46),
			data_in            => s_data_in(14,46),
			data_out           => s_data_out(14,46),
			out1               => s_out1(14,46),
			out2               => s_out2(14,46),
			lock_lower_row_out => s_locks_lower_out(14,46),
			lock_lower_row_in  => s_locks_lower_in(14,46),
			in1                => s_in1(14,46),
			in2                => s_in2(14,46),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(46)
		);
	s_in1(14,46)            <= s_out1(15,46);
	s_in2(14,46)            <= s_out2(15,47);
	s_locks_lower_in(14,46) <= s_locks_lower_out(15,46);

		normal_cell_14_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,47),
			fetch              => s_fetch(14,47),
			data_in            => s_data_in(14,47),
			data_out           => s_data_out(14,47),
			out1               => s_out1(14,47),
			out2               => s_out2(14,47),
			lock_lower_row_out => s_locks_lower_out(14,47),
			lock_lower_row_in  => s_locks_lower_in(14,47),
			in1                => s_in1(14,47),
			in2                => s_in2(14,47),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(47)
		);
	s_in1(14,47)            <= s_out1(15,47);
	s_in2(14,47)            <= s_out2(15,48);
	s_locks_lower_in(14,47) <= s_locks_lower_out(15,47);

		normal_cell_14_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,48),
			fetch              => s_fetch(14,48),
			data_in            => s_data_in(14,48),
			data_out           => s_data_out(14,48),
			out1               => s_out1(14,48),
			out2               => s_out2(14,48),
			lock_lower_row_out => s_locks_lower_out(14,48),
			lock_lower_row_in  => s_locks_lower_in(14,48),
			in1                => s_in1(14,48),
			in2                => s_in2(14,48),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(48)
		);
	s_in1(14,48)            <= s_out1(15,48);
	s_in2(14,48)            <= s_out2(15,49);
	s_locks_lower_in(14,48) <= s_locks_lower_out(15,48);

		normal_cell_14_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,49),
			fetch              => s_fetch(14,49),
			data_in            => s_data_in(14,49),
			data_out           => s_data_out(14,49),
			out1               => s_out1(14,49),
			out2               => s_out2(14,49),
			lock_lower_row_out => s_locks_lower_out(14,49),
			lock_lower_row_in  => s_locks_lower_in(14,49),
			in1                => s_in1(14,49),
			in2                => s_in2(14,49),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(49)
		);
	s_in1(14,49)            <= s_out1(15,49);
	s_in2(14,49)            <= s_out2(15,50);
	s_locks_lower_in(14,49) <= s_locks_lower_out(15,49);

		normal_cell_14_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,50),
			fetch              => s_fetch(14,50),
			data_in            => s_data_in(14,50),
			data_out           => s_data_out(14,50),
			out1               => s_out1(14,50),
			out2               => s_out2(14,50),
			lock_lower_row_out => s_locks_lower_out(14,50),
			lock_lower_row_in  => s_locks_lower_in(14,50),
			in1                => s_in1(14,50),
			in2                => s_in2(14,50),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(50)
		);
	s_in1(14,50)            <= s_out1(15,50);
	s_in2(14,50)            <= s_out2(15,51);
	s_locks_lower_in(14,50) <= s_locks_lower_out(15,50);

		normal_cell_14_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,51),
			fetch              => s_fetch(14,51),
			data_in            => s_data_in(14,51),
			data_out           => s_data_out(14,51),
			out1               => s_out1(14,51),
			out2               => s_out2(14,51),
			lock_lower_row_out => s_locks_lower_out(14,51),
			lock_lower_row_in  => s_locks_lower_in(14,51),
			in1                => s_in1(14,51),
			in2                => s_in2(14,51),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(51)
		);
	s_in1(14,51)            <= s_out1(15,51);
	s_in2(14,51)            <= s_out2(15,52);
	s_locks_lower_in(14,51) <= s_locks_lower_out(15,51);

		normal_cell_14_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,52),
			fetch              => s_fetch(14,52),
			data_in            => s_data_in(14,52),
			data_out           => s_data_out(14,52),
			out1               => s_out1(14,52),
			out2               => s_out2(14,52),
			lock_lower_row_out => s_locks_lower_out(14,52),
			lock_lower_row_in  => s_locks_lower_in(14,52),
			in1                => s_in1(14,52),
			in2                => s_in2(14,52),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(52)
		);
	s_in1(14,52)            <= s_out1(15,52);
	s_in2(14,52)            <= s_out2(15,53);
	s_locks_lower_in(14,52) <= s_locks_lower_out(15,52);

		normal_cell_14_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,53),
			fetch              => s_fetch(14,53),
			data_in            => s_data_in(14,53),
			data_out           => s_data_out(14,53),
			out1               => s_out1(14,53),
			out2               => s_out2(14,53),
			lock_lower_row_out => s_locks_lower_out(14,53),
			lock_lower_row_in  => s_locks_lower_in(14,53),
			in1                => s_in1(14,53),
			in2                => s_in2(14,53),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(53)
		);
	s_in1(14,53)            <= s_out1(15,53);
	s_in2(14,53)            <= s_out2(15,54);
	s_locks_lower_in(14,53) <= s_locks_lower_out(15,53);

		normal_cell_14_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,54),
			fetch              => s_fetch(14,54),
			data_in            => s_data_in(14,54),
			data_out           => s_data_out(14,54),
			out1               => s_out1(14,54),
			out2               => s_out2(14,54),
			lock_lower_row_out => s_locks_lower_out(14,54),
			lock_lower_row_in  => s_locks_lower_in(14,54),
			in1                => s_in1(14,54),
			in2                => s_in2(14,54),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(54)
		);
	s_in1(14,54)            <= s_out1(15,54);
	s_in2(14,54)            <= s_out2(15,55);
	s_locks_lower_in(14,54) <= s_locks_lower_out(15,54);

		normal_cell_14_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,55),
			fetch              => s_fetch(14,55),
			data_in            => s_data_in(14,55),
			data_out           => s_data_out(14,55),
			out1               => s_out1(14,55),
			out2               => s_out2(14,55),
			lock_lower_row_out => s_locks_lower_out(14,55),
			lock_lower_row_in  => s_locks_lower_in(14,55),
			in1                => s_in1(14,55),
			in2                => s_in2(14,55),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(55)
		);
	s_in1(14,55)            <= s_out1(15,55);
	s_in2(14,55)            <= s_out2(15,56);
	s_locks_lower_in(14,55) <= s_locks_lower_out(15,55);

		normal_cell_14_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,56),
			fetch              => s_fetch(14,56),
			data_in            => s_data_in(14,56),
			data_out           => s_data_out(14,56),
			out1               => s_out1(14,56),
			out2               => s_out2(14,56),
			lock_lower_row_out => s_locks_lower_out(14,56),
			lock_lower_row_in  => s_locks_lower_in(14,56),
			in1                => s_in1(14,56),
			in2                => s_in2(14,56),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(56)
		);
	s_in1(14,56)            <= s_out1(15,56);
	s_in2(14,56)            <= s_out2(15,57);
	s_locks_lower_in(14,56) <= s_locks_lower_out(15,56);

		normal_cell_14_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,57),
			fetch              => s_fetch(14,57),
			data_in            => s_data_in(14,57),
			data_out           => s_data_out(14,57),
			out1               => s_out1(14,57),
			out2               => s_out2(14,57),
			lock_lower_row_out => s_locks_lower_out(14,57),
			lock_lower_row_in  => s_locks_lower_in(14,57),
			in1                => s_in1(14,57),
			in2                => s_in2(14,57),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(57)
		);
	s_in1(14,57)            <= s_out1(15,57);
	s_in2(14,57)            <= s_out2(15,58);
	s_locks_lower_in(14,57) <= s_locks_lower_out(15,57);

		normal_cell_14_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,58),
			fetch              => s_fetch(14,58),
			data_in            => s_data_in(14,58),
			data_out           => s_data_out(14,58),
			out1               => s_out1(14,58),
			out2               => s_out2(14,58),
			lock_lower_row_out => s_locks_lower_out(14,58),
			lock_lower_row_in  => s_locks_lower_in(14,58),
			in1                => s_in1(14,58),
			in2                => s_in2(14,58),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(58)
		);
	s_in1(14,58)            <= s_out1(15,58);
	s_in2(14,58)            <= s_out2(15,59);
	s_locks_lower_in(14,58) <= s_locks_lower_out(15,58);

		normal_cell_14_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,59),
			fetch              => s_fetch(14,59),
			data_in            => s_data_in(14,59),
			data_out           => s_data_out(14,59),
			out1               => s_out1(14,59),
			out2               => s_out2(14,59),
			lock_lower_row_out => s_locks_lower_out(14,59),
			lock_lower_row_in  => s_locks_lower_in(14,59),
			in1                => s_in1(14,59),
			in2                => s_in2(14,59),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(59)
		);
	s_in1(14,59)            <= s_out1(15,59);
	s_in2(14,59)            <= s_out2(15,60);
	s_locks_lower_in(14,59) <= s_locks_lower_out(15,59);

		last_col_cell_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(14,60),
			fetch              => s_fetch(14,60),
			data_in            => s_data_in(14,60),
			data_out           => s_data_out(14,60),
			out1               => s_out1(14,60),
			out2               => s_out2(14,60),
			lock_lower_row_out => s_locks_lower_out(14,60),
			lock_lower_row_in  => s_locks_lower_in(14,60),
			in1                => s_in1(14,60),
			in2                => (others => '0'),
			lock_row           => s_locks(14),
			piv_found          => s_piv_found,
			row_data           => s_row_data(14),
			col_data           => s_col_data(60)
		);
	s_in1(14,60)            <= s_out1(15,60);
	s_locks_lower_in(14,60) <= s_locks_lower_out(15,60);

		normal_cell_15_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,1),
			fetch              => s_fetch(15,1),
			data_in            => s_data_in(15,1),
			data_out           => s_data_out(15,1),
			out1               => s_out1(15,1),
			out2               => s_out2(15,1),
			lock_lower_row_out => s_locks_lower_out(15,1),
			lock_lower_row_in  => s_locks_lower_in(15,1),
			in1                => s_in1(15,1),
			in2                => s_in2(15,1),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(1)
		);
	s_in1(15,1)            <= s_out1(16,1);
	s_in2(15,1)            <= s_out2(16,2);
	s_locks_lower_in(15,1) <= s_locks_lower_out(16,1);

		normal_cell_15_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,2),
			fetch              => s_fetch(15,2),
			data_in            => s_data_in(15,2),
			data_out           => s_data_out(15,2),
			out1               => s_out1(15,2),
			out2               => s_out2(15,2),
			lock_lower_row_out => s_locks_lower_out(15,2),
			lock_lower_row_in  => s_locks_lower_in(15,2),
			in1                => s_in1(15,2),
			in2                => s_in2(15,2),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(2)
		);
	s_in1(15,2)            <= s_out1(16,2);
	s_in2(15,2)            <= s_out2(16,3);
	s_locks_lower_in(15,2) <= s_locks_lower_out(16,2);

		normal_cell_15_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,3),
			fetch              => s_fetch(15,3),
			data_in            => s_data_in(15,3),
			data_out           => s_data_out(15,3),
			out1               => s_out1(15,3),
			out2               => s_out2(15,3),
			lock_lower_row_out => s_locks_lower_out(15,3),
			lock_lower_row_in  => s_locks_lower_in(15,3),
			in1                => s_in1(15,3),
			in2                => s_in2(15,3),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(3)
		);
	s_in1(15,3)            <= s_out1(16,3);
	s_in2(15,3)            <= s_out2(16,4);
	s_locks_lower_in(15,3) <= s_locks_lower_out(16,3);

		normal_cell_15_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,4),
			fetch              => s_fetch(15,4),
			data_in            => s_data_in(15,4),
			data_out           => s_data_out(15,4),
			out1               => s_out1(15,4),
			out2               => s_out2(15,4),
			lock_lower_row_out => s_locks_lower_out(15,4),
			lock_lower_row_in  => s_locks_lower_in(15,4),
			in1                => s_in1(15,4),
			in2                => s_in2(15,4),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(4)
		);
	s_in1(15,4)            <= s_out1(16,4);
	s_in2(15,4)            <= s_out2(16,5);
	s_locks_lower_in(15,4) <= s_locks_lower_out(16,4);

		normal_cell_15_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,5),
			fetch              => s_fetch(15,5),
			data_in            => s_data_in(15,5),
			data_out           => s_data_out(15,5),
			out1               => s_out1(15,5),
			out2               => s_out2(15,5),
			lock_lower_row_out => s_locks_lower_out(15,5),
			lock_lower_row_in  => s_locks_lower_in(15,5),
			in1                => s_in1(15,5),
			in2                => s_in2(15,5),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(5)
		);
	s_in1(15,5)            <= s_out1(16,5);
	s_in2(15,5)            <= s_out2(16,6);
	s_locks_lower_in(15,5) <= s_locks_lower_out(16,5);

		normal_cell_15_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,6),
			fetch              => s_fetch(15,6),
			data_in            => s_data_in(15,6),
			data_out           => s_data_out(15,6),
			out1               => s_out1(15,6),
			out2               => s_out2(15,6),
			lock_lower_row_out => s_locks_lower_out(15,6),
			lock_lower_row_in  => s_locks_lower_in(15,6),
			in1                => s_in1(15,6),
			in2                => s_in2(15,6),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(6)
		);
	s_in1(15,6)            <= s_out1(16,6);
	s_in2(15,6)            <= s_out2(16,7);
	s_locks_lower_in(15,6) <= s_locks_lower_out(16,6);

		normal_cell_15_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,7),
			fetch              => s_fetch(15,7),
			data_in            => s_data_in(15,7),
			data_out           => s_data_out(15,7),
			out1               => s_out1(15,7),
			out2               => s_out2(15,7),
			lock_lower_row_out => s_locks_lower_out(15,7),
			lock_lower_row_in  => s_locks_lower_in(15,7),
			in1                => s_in1(15,7),
			in2                => s_in2(15,7),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(7)
		);
	s_in1(15,7)            <= s_out1(16,7);
	s_in2(15,7)            <= s_out2(16,8);
	s_locks_lower_in(15,7) <= s_locks_lower_out(16,7);

		normal_cell_15_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,8),
			fetch              => s_fetch(15,8),
			data_in            => s_data_in(15,8),
			data_out           => s_data_out(15,8),
			out1               => s_out1(15,8),
			out2               => s_out2(15,8),
			lock_lower_row_out => s_locks_lower_out(15,8),
			lock_lower_row_in  => s_locks_lower_in(15,8),
			in1                => s_in1(15,8),
			in2                => s_in2(15,8),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(8)
		);
	s_in1(15,8)            <= s_out1(16,8);
	s_in2(15,8)            <= s_out2(16,9);
	s_locks_lower_in(15,8) <= s_locks_lower_out(16,8);

		normal_cell_15_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,9),
			fetch              => s_fetch(15,9),
			data_in            => s_data_in(15,9),
			data_out           => s_data_out(15,9),
			out1               => s_out1(15,9),
			out2               => s_out2(15,9),
			lock_lower_row_out => s_locks_lower_out(15,9),
			lock_lower_row_in  => s_locks_lower_in(15,9),
			in1                => s_in1(15,9),
			in2                => s_in2(15,9),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(9)
		);
	s_in1(15,9)            <= s_out1(16,9);
	s_in2(15,9)            <= s_out2(16,10);
	s_locks_lower_in(15,9) <= s_locks_lower_out(16,9);

		normal_cell_15_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,10),
			fetch              => s_fetch(15,10),
			data_in            => s_data_in(15,10),
			data_out           => s_data_out(15,10),
			out1               => s_out1(15,10),
			out2               => s_out2(15,10),
			lock_lower_row_out => s_locks_lower_out(15,10),
			lock_lower_row_in  => s_locks_lower_in(15,10),
			in1                => s_in1(15,10),
			in2                => s_in2(15,10),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(10)
		);
	s_in1(15,10)            <= s_out1(16,10);
	s_in2(15,10)            <= s_out2(16,11);
	s_locks_lower_in(15,10) <= s_locks_lower_out(16,10);

		normal_cell_15_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,11),
			fetch              => s_fetch(15,11),
			data_in            => s_data_in(15,11),
			data_out           => s_data_out(15,11),
			out1               => s_out1(15,11),
			out2               => s_out2(15,11),
			lock_lower_row_out => s_locks_lower_out(15,11),
			lock_lower_row_in  => s_locks_lower_in(15,11),
			in1                => s_in1(15,11),
			in2                => s_in2(15,11),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(11)
		);
	s_in1(15,11)            <= s_out1(16,11);
	s_in2(15,11)            <= s_out2(16,12);
	s_locks_lower_in(15,11) <= s_locks_lower_out(16,11);

		normal_cell_15_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,12),
			fetch              => s_fetch(15,12),
			data_in            => s_data_in(15,12),
			data_out           => s_data_out(15,12),
			out1               => s_out1(15,12),
			out2               => s_out2(15,12),
			lock_lower_row_out => s_locks_lower_out(15,12),
			lock_lower_row_in  => s_locks_lower_in(15,12),
			in1                => s_in1(15,12),
			in2                => s_in2(15,12),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(12)
		);
	s_in1(15,12)            <= s_out1(16,12);
	s_in2(15,12)            <= s_out2(16,13);
	s_locks_lower_in(15,12) <= s_locks_lower_out(16,12);

		normal_cell_15_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,13),
			fetch              => s_fetch(15,13),
			data_in            => s_data_in(15,13),
			data_out           => s_data_out(15,13),
			out1               => s_out1(15,13),
			out2               => s_out2(15,13),
			lock_lower_row_out => s_locks_lower_out(15,13),
			lock_lower_row_in  => s_locks_lower_in(15,13),
			in1                => s_in1(15,13),
			in2                => s_in2(15,13),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(13)
		);
	s_in1(15,13)            <= s_out1(16,13);
	s_in2(15,13)            <= s_out2(16,14);
	s_locks_lower_in(15,13) <= s_locks_lower_out(16,13);

		normal_cell_15_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,14),
			fetch              => s_fetch(15,14),
			data_in            => s_data_in(15,14),
			data_out           => s_data_out(15,14),
			out1               => s_out1(15,14),
			out2               => s_out2(15,14),
			lock_lower_row_out => s_locks_lower_out(15,14),
			lock_lower_row_in  => s_locks_lower_in(15,14),
			in1                => s_in1(15,14),
			in2                => s_in2(15,14),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(14)
		);
	s_in1(15,14)            <= s_out1(16,14);
	s_in2(15,14)            <= s_out2(16,15);
	s_locks_lower_in(15,14) <= s_locks_lower_out(16,14);

		normal_cell_15_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,15),
			fetch              => s_fetch(15,15),
			data_in            => s_data_in(15,15),
			data_out           => s_data_out(15,15),
			out1               => s_out1(15,15),
			out2               => s_out2(15,15),
			lock_lower_row_out => s_locks_lower_out(15,15),
			lock_lower_row_in  => s_locks_lower_in(15,15),
			in1                => s_in1(15,15),
			in2                => s_in2(15,15),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(15)
		);
	s_in1(15,15)            <= s_out1(16,15);
	s_in2(15,15)            <= s_out2(16,16);
	s_locks_lower_in(15,15) <= s_locks_lower_out(16,15);

		normal_cell_15_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,16),
			fetch              => s_fetch(15,16),
			data_in            => s_data_in(15,16),
			data_out           => s_data_out(15,16),
			out1               => s_out1(15,16),
			out2               => s_out2(15,16),
			lock_lower_row_out => s_locks_lower_out(15,16),
			lock_lower_row_in  => s_locks_lower_in(15,16),
			in1                => s_in1(15,16),
			in2                => s_in2(15,16),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(16)
		);
	s_in1(15,16)            <= s_out1(16,16);
	s_in2(15,16)            <= s_out2(16,17);
	s_locks_lower_in(15,16) <= s_locks_lower_out(16,16);

		normal_cell_15_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,17),
			fetch              => s_fetch(15,17),
			data_in            => s_data_in(15,17),
			data_out           => s_data_out(15,17),
			out1               => s_out1(15,17),
			out2               => s_out2(15,17),
			lock_lower_row_out => s_locks_lower_out(15,17),
			lock_lower_row_in  => s_locks_lower_in(15,17),
			in1                => s_in1(15,17),
			in2                => s_in2(15,17),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(17)
		);
	s_in1(15,17)            <= s_out1(16,17);
	s_in2(15,17)            <= s_out2(16,18);
	s_locks_lower_in(15,17) <= s_locks_lower_out(16,17);

		normal_cell_15_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,18),
			fetch              => s_fetch(15,18),
			data_in            => s_data_in(15,18),
			data_out           => s_data_out(15,18),
			out1               => s_out1(15,18),
			out2               => s_out2(15,18),
			lock_lower_row_out => s_locks_lower_out(15,18),
			lock_lower_row_in  => s_locks_lower_in(15,18),
			in1                => s_in1(15,18),
			in2                => s_in2(15,18),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(18)
		);
	s_in1(15,18)            <= s_out1(16,18);
	s_in2(15,18)            <= s_out2(16,19);
	s_locks_lower_in(15,18) <= s_locks_lower_out(16,18);

		normal_cell_15_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,19),
			fetch              => s_fetch(15,19),
			data_in            => s_data_in(15,19),
			data_out           => s_data_out(15,19),
			out1               => s_out1(15,19),
			out2               => s_out2(15,19),
			lock_lower_row_out => s_locks_lower_out(15,19),
			lock_lower_row_in  => s_locks_lower_in(15,19),
			in1                => s_in1(15,19),
			in2                => s_in2(15,19),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(19)
		);
	s_in1(15,19)            <= s_out1(16,19);
	s_in2(15,19)            <= s_out2(16,20);
	s_locks_lower_in(15,19) <= s_locks_lower_out(16,19);

		normal_cell_15_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,20),
			fetch              => s_fetch(15,20),
			data_in            => s_data_in(15,20),
			data_out           => s_data_out(15,20),
			out1               => s_out1(15,20),
			out2               => s_out2(15,20),
			lock_lower_row_out => s_locks_lower_out(15,20),
			lock_lower_row_in  => s_locks_lower_in(15,20),
			in1                => s_in1(15,20),
			in2                => s_in2(15,20),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(20)
		);
	s_in1(15,20)            <= s_out1(16,20);
	s_in2(15,20)            <= s_out2(16,21);
	s_locks_lower_in(15,20) <= s_locks_lower_out(16,20);

		normal_cell_15_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,21),
			fetch              => s_fetch(15,21),
			data_in            => s_data_in(15,21),
			data_out           => s_data_out(15,21),
			out1               => s_out1(15,21),
			out2               => s_out2(15,21),
			lock_lower_row_out => s_locks_lower_out(15,21),
			lock_lower_row_in  => s_locks_lower_in(15,21),
			in1                => s_in1(15,21),
			in2                => s_in2(15,21),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(21)
		);
	s_in1(15,21)            <= s_out1(16,21);
	s_in2(15,21)            <= s_out2(16,22);
	s_locks_lower_in(15,21) <= s_locks_lower_out(16,21);

		normal_cell_15_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,22),
			fetch              => s_fetch(15,22),
			data_in            => s_data_in(15,22),
			data_out           => s_data_out(15,22),
			out1               => s_out1(15,22),
			out2               => s_out2(15,22),
			lock_lower_row_out => s_locks_lower_out(15,22),
			lock_lower_row_in  => s_locks_lower_in(15,22),
			in1                => s_in1(15,22),
			in2                => s_in2(15,22),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(22)
		);
	s_in1(15,22)            <= s_out1(16,22);
	s_in2(15,22)            <= s_out2(16,23);
	s_locks_lower_in(15,22) <= s_locks_lower_out(16,22);

		normal_cell_15_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,23),
			fetch              => s_fetch(15,23),
			data_in            => s_data_in(15,23),
			data_out           => s_data_out(15,23),
			out1               => s_out1(15,23),
			out2               => s_out2(15,23),
			lock_lower_row_out => s_locks_lower_out(15,23),
			lock_lower_row_in  => s_locks_lower_in(15,23),
			in1                => s_in1(15,23),
			in2                => s_in2(15,23),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(23)
		);
	s_in1(15,23)            <= s_out1(16,23);
	s_in2(15,23)            <= s_out2(16,24);
	s_locks_lower_in(15,23) <= s_locks_lower_out(16,23);

		normal_cell_15_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,24),
			fetch              => s_fetch(15,24),
			data_in            => s_data_in(15,24),
			data_out           => s_data_out(15,24),
			out1               => s_out1(15,24),
			out2               => s_out2(15,24),
			lock_lower_row_out => s_locks_lower_out(15,24),
			lock_lower_row_in  => s_locks_lower_in(15,24),
			in1                => s_in1(15,24),
			in2                => s_in2(15,24),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(24)
		);
	s_in1(15,24)            <= s_out1(16,24);
	s_in2(15,24)            <= s_out2(16,25);
	s_locks_lower_in(15,24) <= s_locks_lower_out(16,24);

		normal_cell_15_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,25),
			fetch              => s_fetch(15,25),
			data_in            => s_data_in(15,25),
			data_out           => s_data_out(15,25),
			out1               => s_out1(15,25),
			out2               => s_out2(15,25),
			lock_lower_row_out => s_locks_lower_out(15,25),
			lock_lower_row_in  => s_locks_lower_in(15,25),
			in1                => s_in1(15,25),
			in2                => s_in2(15,25),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(25)
		);
	s_in1(15,25)            <= s_out1(16,25);
	s_in2(15,25)            <= s_out2(16,26);
	s_locks_lower_in(15,25) <= s_locks_lower_out(16,25);

		normal_cell_15_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,26),
			fetch              => s_fetch(15,26),
			data_in            => s_data_in(15,26),
			data_out           => s_data_out(15,26),
			out1               => s_out1(15,26),
			out2               => s_out2(15,26),
			lock_lower_row_out => s_locks_lower_out(15,26),
			lock_lower_row_in  => s_locks_lower_in(15,26),
			in1                => s_in1(15,26),
			in2                => s_in2(15,26),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(26)
		);
	s_in1(15,26)            <= s_out1(16,26);
	s_in2(15,26)            <= s_out2(16,27);
	s_locks_lower_in(15,26) <= s_locks_lower_out(16,26);

		normal_cell_15_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,27),
			fetch              => s_fetch(15,27),
			data_in            => s_data_in(15,27),
			data_out           => s_data_out(15,27),
			out1               => s_out1(15,27),
			out2               => s_out2(15,27),
			lock_lower_row_out => s_locks_lower_out(15,27),
			lock_lower_row_in  => s_locks_lower_in(15,27),
			in1                => s_in1(15,27),
			in2                => s_in2(15,27),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(27)
		);
	s_in1(15,27)            <= s_out1(16,27);
	s_in2(15,27)            <= s_out2(16,28);
	s_locks_lower_in(15,27) <= s_locks_lower_out(16,27);

		normal_cell_15_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,28),
			fetch              => s_fetch(15,28),
			data_in            => s_data_in(15,28),
			data_out           => s_data_out(15,28),
			out1               => s_out1(15,28),
			out2               => s_out2(15,28),
			lock_lower_row_out => s_locks_lower_out(15,28),
			lock_lower_row_in  => s_locks_lower_in(15,28),
			in1                => s_in1(15,28),
			in2                => s_in2(15,28),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(28)
		);
	s_in1(15,28)            <= s_out1(16,28);
	s_in2(15,28)            <= s_out2(16,29);
	s_locks_lower_in(15,28) <= s_locks_lower_out(16,28);

		normal_cell_15_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,29),
			fetch              => s_fetch(15,29),
			data_in            => s_data_in(15,29),
			data_out           => s_data_out(15,29),
			out1               => s_out1(15,29),
			out2               => s_out2(15,29),
			lock_lower_row_out => s_locks_lower_out(15,29),
			lock_lower_row_in  => s_locks_lower_in(15,29),
			in1                => s_in1(15,29),
			in2                => s_in2(15,29),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(29)
		);
	s_in1(15,29)            <= s_out1(16,29);
	s_in2(15,29)            <= s_out2(16,30);
	s_locks_lower_in(15,29) <= s_locks_lower_out(16,29);

		normal_cell_15_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,30),
			fetch              => s_fetch(15,30),
			data_in            => s_data_in(15,30),
			data_out           => s_data_out(15,30),
			out1               => s_out1(15,30),
			out2               => s_out2(15,30),
			lock_lower_row_out => s_locks_lower_out(15,30),
			lock_lower_row_in  => s_locks_lower_in(15,30),
			in1                => s_in1(15,30),
			in2                => s_in2(15,30),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(30)
		);
	s_in1(15,30)            <= s_out1(16,30);
	s_in2(15,30)            <= s_out2(16,31);
	s_locks_lower_in(15,30) <= s_locks_lower_out(16,30);

		normal_cell_15_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,31),
			fetch              => s_fetch(15,31),
			data_in            => s_data_in(15,31),
			data_out           => s_data_out(15,31),
			out1               => s_out1(15,31),
			out2               => s_out2(15,31),
			lock_lower_row_out => s_locks_lower_out(15,31),
			lock_lower_row_in  => s_locks_lower_in(15,31),
			in1                => s_in1(15,31),
			in2                => s_in2(15,31),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(31)
		);
	s_in1(15,31)            <= s_out1(16,31);
	s_in2(15,31)            <= s_out2(16,32);
	s_locks_lower_in(15,31) <= s_locks_lower_out(16,31);

		normal_cell_15_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,32),
			fetch              => s_fetch(15,32),
			data_in            => s_data_in(15,32),
			data_out           => s_data_out(15,32),
			out1               => s_out1(15,32),
			out2               => s_out2(15,32),
			lock_lower_row_out => s_locks_lower_out(15,32),
			lock_lower_row_in  => s_locks_lower_in(15,32),
			in1                => s_in1(15,32),
			in2                => s_in2(15,32),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(32)
		);
	s_in1(15,32)            <= s_out1(16,32);
	s_in2(15,32)            <= s_out2(16,33);
	s_locks_lower_in(15,32) <= s_locks_lower_out(16,32);

		normal_cell_15_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,33),
			fetch              => s_fetch(15,33),
			data_in            => s_data_in(15,33),
			data_out           => s_data_out(15,33),
			out1               => s_out1(15,33),
			out2               => s_out2(15,33),
			lock_lower_row_out => s_locks_lower_out(15,33),
			lock_lower_row_in  => s_locks_lower_in(15,33),
			in1                => s_in1(15,33),
			in2                => s_in2(15,33),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(33)
		);
	s_in1(15,33)            <= s_out1(16,33);
	s_in2(15,33)            <= s_out2(16,34);
	s_locks_lower_in(15,33) <= s_locks_lower_out(16,33);

		normal_cell_15_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,34),
			fetch              => s_fetch(15,34),
			data_in            => s_data_in(15,34),
			data_out           => s_data_out(15,34),
			out1               => s_out1(15,34),
			out2               => s_out2(15,34),
			lock_lower_row_out => s_locks_lower_out(15,34),
			lock_lower_row_in  => s_locks_lower_in(15,34),
			in1                => s_in1(15,34),
			in2                => s_in2(15,34),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(34)
		);
	s_in1(15,34)            <= s_out1(16,34);
	s_in2(15,34)            <= s_out2(16,35);
	s_locks_lower_in(15,34) <= s_locks_lower_out(16,34);

		normal_cell_15_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,35),
			fetch              => s_fetch(15,35),
			data_in            => s_data_in(15,35),
			data_out           => s_data_out(15,35),
			out1               => s_out1(15,35),
			out2               => s_out2(15,35),
			lock_lower_row_out => s_locks_lower_out(15,35),
			lock_lower_row_in  => s_locks_lower_in(15,35),
			in1                => s_in1(15,35),
			in2                => s_in2(15,35),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(35)
		);
	s_in1(15,35)            <= s_out1(16,35);
	s_in2(15,35)            <= s_out2(16,36);
	s_locks_lower_in(15,35) <= s_locks_lower_out(16,35);

		normal_cell_15_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,36),
			fetch              => s_fetch(15,36),
			data_in            => s_data_in(15,36),
			data_out           => s_data_out(15,36),
			out1               => s_out1(15,36),
			out2               => s_out2(15,36),
			lock_lower_row_out => s_locks_lower_out(15,36),
			lock_lower_row_in  => s_locks_lower_in(15,36),
			in1                => s_in1(15,36),
			in2                => s_in2(15,36),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(36)
		);
	s_in1(15,36)            <= s_out1(16,36);
	s_in2(15,36)            <= s_out2(16,37);
	s_locks_lower_in(15,36) <= s_locks_lower_out(16,36);

		normal_cell_15_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,37),
			fetch              => s_fetch(15,37),
			data_in            => s_data_in(15,37),
			data_out           => s_data_out(15,37),
			out1               => s_out1(15,37),
			out2               => s_out2(15,37),
			lock_lower_row_out => s_locks_lower_out(15,37),
			lock_lower_row_in  => s_locks_lower_in(15,37),
			in1                => s_in1(15,37),
			in2                => s_in2(15,37),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(37)
		);
	s_in1(15,37)            <= s_out1(16,37);
	s_in2(15,37)            <= s_out2(16,38);
	s_locks_lower_in(15,37) <= s_locks_lower_out(16,37);

		normal_cell_15_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,38),
			fetch              => s_fetch(15,38),
			data_in            => s_data_in(15,38),
			data_out           => s_data_out(15,38),
			out1               => s_out1(15,38),
			out2               => s_out2(15,38),
			lock_lower_row_out => s_locks_lower_out(15,38),
			lock_lower_row_in  => s_locks_lower_in(15,38),
			in1                => s_in1(15,38),
			in2                => s_in2(15,38),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(38)
		);
	s_in1(15,38)            <= s_out1(16,38);
	s_in2(15,38)            <= s_out2(16,39);
	s_locks_lower_in(15,38) <= s_locks_lower_out(16,38);

		normal_cell_15_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,39),
			fetch              => s_fetch(15,39),
			data_in            => s_data_in(15,39),
			data_out           => s_data_out(15,39),
			out1               => s_out1(15,39),
			out2               => s_out2(15,39),
			lock_lower_row_out => s_locks_lower_out(15,39),
			lock_lower_row_in  => s_locks_lower_in(15,39),
			in1                => s_in1(15,39),
			in2                => s_in2(15,39),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(39)
		);
	s_in1(15,39)            <= s_out1(16,39);
	s_in2(15,39)            <= s_out2(16,40);
	s_locks_lower_in(15,39) <= s_locks_lower_out(16,39);

		normal_cell_15_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,40),
			fetch              => s_fetch(15,40),
			data_in            => s_data_in(15,40),
			data_out           => s_data_out(15,40),
			out1               => s_out1(15,40),
			out2               => s_out2(15,40),
			lock_lower_row_out => s_locks_lower_out(15,40),
			lock_lower_row_in  => s_locks_lower_in(15,40),
			in1                => s_in1(15,40),
			in2                => s_in2(15,40),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(40)
		);
	s_in1(15,40)            <= s_out1(16,40);
	s_in2(15,40)            <= s_out2(16,41);
	s_locks_lower_in(15,40) <= s_locks_lower_out(16,40);

		normal_cell_15_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,41),
			fetch              => s_fetch(15,41),
			data_in            => s_data_in(15,41),
			data_out           => s_data_out(15,41),
			out1               => s_out1(15,41),
			out2               => s_out2(15,41),
			lock_lower_row_out => s_locks_lower_out(15,41),
			lock_lower_row_in  => s_locks_lower_in(15,41),
			in1                => s_in1(15,41),
			in2                => s_in2(15,41),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(41)
		);
	s_in1(15,41)            <= s_out1(16,41);
	s_in2(15,41)            <= s_out2(16,42);
	s_locks_lower_in(15,41) <= s_locks_lower_out(16,41);

		normal_cell_15_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,42),
			fetch              => s_fetch(15,42),
			data_in            => s_data_in(15,42),
			data_out           => s_data_out(15,42),
			out1               => s_out1(15,42),
			out2               => s_out2(15,42),
			lock_lower_row_out => s_locks_lower_out(15,42),
			lock_lower_row_in  => s_locks_lower_in(15,42),
			in1                => s_in1(15,42),
			in2                => s_in2(15,42),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(42)
		);
	s_in1(15,42)            <= s_out1(16,42);
	s_in2(15,42)            <= s_out2(16,43);
	s_locks_lower_in(15,42) <= s_locks_lower_out(16,42);

		normal_cell_15_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,43),
			fetch              => s_fetch(15,43),
			data_in            => s_data_in(15,43),
			data_out           => s_data_out(15,43),
			out1               => s_out1(15,43),
			out2               => s_out2(15,43),
			lock_lower_row_out => s_locks_lower_out(15,43),
			lock_lower_row_in  => s_locks_lower_in(15,43),
			in1                => s_in1(15,43),
			in2                => s_in2(15,43),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(43)
		);
	s_in1(15,43)            <= s_out1(16,43);
	s_in2(15,43)            <= s_out2(16,44);
	s_locks_lower_in(15,43) <= s_locks_lower_out(16,43);

		normal_cell_15_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,44),
			fetch              => s_fetch(15,44),
			data_in            => s_data_in(15,44),
			data_out           => s_data_out(15,44),
			out1               => s_out1(15,44),
			out2               => s_out2(15,44),
			lock_lower_row_out => s_locks_lower_out(15,44),
			lock_lower_row_in  => s_locks_lower_in(15,44),
			in1                => s_in1(15,44),
			in2                => s_in2(15,44),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(44)
		);
	s_in1(15,44)            <= s_out1(16,44);
	s_in2(15,44)            <= s_out2(16,45);
	s_locks_lower_in(15,44) <= s_locks_lower_out(16,44);

		normal_cell_15_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,45),
			fetch              => s_fetch(15,45),
			data_in            => s_data_in(15,45),
			data_out           => s_data_out(15,45),
			out1               => s_out1(15,45),
			out2               => s_out2(15,45),
			lock_lower_row_out => s_locks_lower_out(15,45),
			lock_lower_row_in  => s_locks_lower_in(15,45),
			in1                => s_in1(15,45),
			in2                => s_in2(15,45),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(45)
		);
	s_in1(15,45)            <= s_out1(16,45);
	s_in2(15,45)            <= s_out2(16,46);
	s_locks_lower_in(15,45) <= s_locks_lower_out(16,45);

		normal_cell_15_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,46),
			fetch              => s_fetch(15,46),
			data_in            => s_data_in(15,46),
			data_out           => s_data_out(15,46),
			out1               => s_out1(15,46),
			out2               => s_out2(15,46),
			lock_lower_row_out => s_locks_lower_out(15,46),
			lock_lower_row_in  => s_locks_lower_in(15,46),
			in1                => s_in1(15,46),
			in2                => s_in2(15,46),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(46)
		);
	s_in1(15,46)            <= s_out1(16,46);
	s_in2(15,46)            <= s_out2(16,47);
	s_locks_lower_in(15,46) <= s_locks_lower_out(16,46);

		normal_cell_15_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,47),
			fetch              => s_fetch(15,47),
			data_in            => s_data_in(15,47),
			data_out           => s_data_out(15,47),
			out1               => s_out1(15,47),
			out2               => s_out2(15,47),
			lock_lower_row_out => s_locks_lower_out(15,47),
			lock_lower_row_in  => s_locks_lower_in(15,47),
			in1                => s_in1(15,47),
			in2                => s_in2(15,47),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(47)
		);
	s_in1(15,47)            <= s_out1(16,47);
	s_in2(15,47)            <= s_out2(16,48);
	s_locks_lower_in(15,47) <= s_locks_lower_out(16,47);

		normal_cell_15_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,48),
			fetch              => s_fetch(15,48),
			data_in            => s_data_in(15,48),
			data_out           => s_data_out(15,48),
			out1               => s_out1(15,48),
			out2               => s_out2(15,48),
			lock_lower_row_out => s_locks_lower_out(15,48),
			lock_lower_row_in  => s_locks_lower_in(15,48),
			in1                => s_in1(15,48),
			in2                => s_in2(15,48),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(48)
		);
	s_in1(15,48)            <= s_out1(16,48);
	s_in2(15,48)            <= s_out2(16,49);
	s_locks_lower_in(15,48) <= s_locks_lower_out(16,48);

		normal_cell_15_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,49),
			fetch              => s_fetch(15,49),
			data_in            => s_data_in(15,49),
			data_out           => s_data_out(15,49),
			out1               => s_out1(15,49),
			out2               => s_out2(15,49),
			lock_lower_row_out => s_locks_lower_out(15,49),
			lock_lower_row_in  => s_locks_lower_in(15,49),
			in1                => s_in1(15,49),
			in2                => s_in2(15,49),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(49)
		);
	s_in1(15,49)            <= s_out1(16,49);
	s_in2(15,49)            <= s_out2(16,50);
	s_locks_lower_in(15,49) <= s_locks_lower_out(16,49);

		normal_cell_15_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,50),
			fetch              => s_fetch(15,50),
			data_in            => s_data_in(15,50),
			data_out           => s_data_out(15,50),
			out1               => s_out1(15,50),
			out2               => s_out2(15,50),
			lock_lower_row_out => s_locks_lower_out(15,50),
			lock_lower_row_in  => s_locks_lower_in(15,50),
			in1                => s_in1(15,50),
			in2                => s_in2(15,50),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(50)
		);
	s_in1(15,50)            <= s_out1(16,50);
	s_in2(15,50)            <= s_out2(16,51);
	s_locks_lower_in(15,50) <= s_locks_lower_out(16,50);

		normal_cell_15_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,51),
			fetch              => s_fetch(15,51),
			data_in            => s_data_in(15,51),
			data_out           => s_data_out(15,51),
			out1               => s_out1(15,51),
			out2               => s_out2(15,51),
			lock_lower_row_out => s_locks_lower_out(15,51),
			lock_lower_row_in  => s_locks_lower_in(15,51),
			in1                => s_in1(15,51),
			in2                => s_in2(15,51),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(51)
		);
	s_in1(15,51)            <= s_out1(16,51);
	s_in2(15,51)            <= s_out2(16,52);
	s_locks_lower_in(15,51) <= s_locks_lower_out(16,51);

		normal_cell_15_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,52),
			fetch              => s_fetch(15,52),
			data_in            => s_data_in(15,52),
			data_out           => s_data_out(15,52),
			out1               => s_out1(15,52),
			out2               => s_out2(15,52),
			lock_lower_row_out => s_locks_lower_out(15,52),
			lock_lower_row_in  => s_locks_lower_in(15,52),
			in1                => s_in1(15,52),
			in2                => s_in2(15,52),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(52)
		);
	s_in1(15,52)            <= s_out1(16,52);
	s_in2(15,52)            <= s_out2(16,53);
	s_locks_lower_in(15,52) <= s_locks_lower_out(16,52);

		normal_cell_15_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,53),
			fetch              => s_fetch(15,53),
			data_in            => s_data_in(15,53),
			data_out           => s_data_out(15,53),
			out1               => s_out1(15,53),
			out2               => s_out2(15,53),
			lock_lower_row_out => s_locks_lower_out(15,53),
			lock_lower_row_in  => s_locks_lower_in(15,53),
			in1                => s_in1(15,53),
			in2                => s_in2(15,53),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(53)
		);
	s_in1(15,53)            <= s_out1(16,53);
	s_in2(15,53)            <= s_out2(16,54);
	s_locks_lower_in(15,53) <= s_locks_lower_out(16,53);

		normal_cell_15_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,54),
			fetch              => s_fetch(15,54),
			data_in            => s_data_in(15,54),
			data_out           => s_data_out(15,54),
			out1               => s_out1(15,54),
			out2               => s_out2(15,54),
			lock_lower_row_out => s_locks_lower_out(15,54),
			lock_lower_row_in  => s_locks_lower_in(15,54),
			in1                => s_in1(15,54),
			in2                => s_in2(15,54),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(54)
		);
	s_in1(15,54)            <= s_out1(16,54);
	s_in2(15,54)            <= s_out2(16,55);
	s_locks_lower_in(15,54) <= s_locks_lower_out(16,54);

		normal_cell_15_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,55),
			fetch              => s_fetch(15,55),
			data_in            => s_data_in(15,55),
			data_out           => s_data_out(15,55),
			out1               => s_out1(15,55),
			out2               => s_out2(15,55),
			lock_lower_row_out => s_locks_lower_out(15,55),
			lock_lower_row_in  => s_locks_lower_in(15,55),
			in1                => s_in1(15,55),
			in2                => s_in2(15,55),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(55)
		);
	s_in1(15,55)            <= s_out1(16,55);
	s_in2(15,55)            <= s_out2(16,56);
	s_locks_lower_in(15,55) <= s_locks_lower_out(16,55);

		normal_cell_15_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,56),
			fetch              => s_fetch(15,56),
			data_in            => s_data_in(15,56),
			data_out           => s_data_out(15,56),
			out1               => s_out1(15,56),
			out2               => s_out2(15,56),
			lock_lower_row_out => s_locks_lower_out(15,56),
			lock_lower_row_in  => s_locks_lower_in(15,56),
			in1                => s_in1(15,56),
			in2                => s_in2(15,56),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(56)
		);
	s_in1(15,56)            <= s_out1(16,56);
	s_in2(15,56)            <= s_out2(16,57);
	s_locks_lower_in(15,56) <= s_locks_lower_out(16,56);

		normal_cell_15_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,57),
			fetch              => s_fetch(15,57),
			data_in            => s_data_in(15,57),
			data_out           => s_data_out(15,57),
			out1               => s_out1(15,57),
			out2               => s_out2(15,57),
			lock_lower_row_out => s_locks_lower_out(15,57),
			lock_lower_row_in  => s_locks_lower_in(15,57),
			in1                => s_in1(15,57),
			in2                => s_in2(15,57),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(57)
		);
	s_in1(15,57)            <= s_out1(16,57);
	s_in2(15,57)            <= s_out2(16,58);
	s_locks_lower_in(15,57) <= s_locks_lower_out(16,57);

		normal_cell_15_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,58),
			fetch              => s_fetch(15,58),
			data_in            => s_data_in(15,58),
			data_out           => s_data_out(15,58),
			out1               => s_out1(15,58),
			out2               => s_out2(15,58),
			lock_lower_row_out => s_locks_lower_out(15,58),
			lock_lower_row_in  => s_locks_lower_in(15,58),
			in1                => s_in1(15,58),
			in2                => s_in2(15,58),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(58)
		);
	s_in1(15,58)            <= s_out1(16,58);
	s_in2(15,58)            <= s_out2(16,59);
	s_locks_lower_in(15,58) <= s_locks_lower_out(16,58);

		normal_cell_15_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,59),
			fetch              => s_fetch(15,59),
			data_in            => s_data_in(15,59),
			data_out           => s_data_out(15,59),
			out1               => s_out1(15,59),
			out2               => s_out2(15,59),
			lock_lower_row_out => s_locks_lower_out(15,59),
			lock_lower_row_in  => s_locks_lower_in(15,59),
			in1                => s_in1(15,59),
			in2                => s_in2(15,59),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(59)
		);
	s_in1(15,59)            <= s_out1(16,59);
	s_in2(15,59)            <= s_out2(16,60);
	s_locks_lower_in(15,59) <= s_locks_lower_out(16,59);

		last_col_cell_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(15,60),
			fetch              => s_fetch(15,60),
			data_in            => s_data_in(15,60),
			data_out           => s_data_out(15,60),
			out1               => s_out1(15,60),
			out2               => s_out2(15,60),
			lock_lower_row_out => s_locks_lower_out(15,60),
			lock_lower_row_in  => s_locks_lower_in(15,60),
			in1                => s_in1(15,60),
			in2                => (others => '0'),
			lock_row           => s_locks(15),
			piv_found          => s_piv_found,
			row_data           => s_row_data(15),
			col_data           => s_col_data(60)
		);
	s_in1(15,60)            <= s_out1(16,60);
	s_locks_lower_in(15,60) <= s_locks_lower_out(16,60);

		normal_cell_16_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,1),
			fetch              => s_fetch(16,1),
			data_in            => s_data_in(16,1),
			data_out           => s_data_out(16,1),
			out1               => s_out1(16,1),
			out2               => s_out2(16,1),
			lock_lower_row_out => s_locks_lower_out(16,1),
			lock_lower_row_in  => s_locks_lower_in(16,1),
			in1                => s_in1(16,1),
			in2                => s_in2(16,1),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(1)
		);
	s_in1(16,1)            <= s_out1(17,1);
	s_in2(16,1)            <= s_out2(17,2);
	s_locks_lower_in(16,1) <= s_locks_lower_out(17,1);

		normal_cell_16_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,2),
			fetch              => s_fetch(16,2),
			data_in            => s_data_in(16,2),
			data_out           => s_data_out(16,2),
			out1               => s_out1(16,2),
			out2               => s_out2(16,2),
			lock_lower_row_out => s_locks_lower_out(16,2),
			lock_lower_row_in  => s_locks_lower_in(16,2),
			in1                => s_in1(16,2),
			in2                => s_in2(16,2),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(2)
		);
	s_in1(16,2)            <= s_out1(17,2);
	s_in2(16,2)            <= s_out2(17,3);
	s_locks_lower_in(16,2) <= s_locks_lower_out(17,2);

		normal_cell_16_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,3),
			fetch              => s_fetch(16,3),
			data_in            => s_data_in(16,3),
			data_out           => s_data_out(16,3),
			out1               => s_out1(16,3),
			out2               => s_out2(16,3),
			lock_lower_row_out => s_locks_lower_out(16,3),
			lock_lower_row_in  => s_locks_lower_in(16,3),
			in1                => s_in1(16,3),
			in2                => s_in2(16,3),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(3)
		);
	s_in1(16,3)            <= s_out1(17,3);
	s_in2(16,3)            <= s_out2(17,4);
	s_locks_lower_in(16,3) <= s_locks_lower_out(17,3);

		normal_cell_16_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,4),
			fetch              => s_fetch(16,4),
			data_in            => s_data_in(16,4),
			data_out           => s_data_out(16,4),
			out1               => s_out1(16,4),
			out2               => s_out2(16,4),
			lock_lower_row_out => s_locks_lower_out(16,4),
			lock_lower_row_in  => s_locks_lower_in(16,4),
			in1                => s_in1(16,4),
			in2                => s_in2(16,4),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(4)
		);
	s_in1(16,4)            <= s_out1(17,4);
	s_in2(16,4)            <= s_out2(17,5);
	s_locks_lower_in(16,4) <= s_locks_lower_out(17,4);

		normal_cell_16_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,5),
			fetch              => s_fetch(16,5),
			data_in            => s_data_in(16,5),
			data_out           => s_data_out(16,5),
			out1               => s_out1(16,5),
			out2               => s_out2(16,5),
			lock_lower_row_out => s_locks_lower_out(16,5),
			lock_lower_row_in  => s_locks_lower_in(16,5),
			in1                => s_in1(16,5),
			in2                => s_in2(16,5),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(5)
		);
	s_in1(16,5)            <= s_out1(17,5);
	s_in2(16,5)            <= s_out2(17,6);
	s_locks_lower_in(16,5) <= s_locks_lower_out(17,5);

		normal_cell_16_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,6),
			fetch              => s_fetch(16,6),
			data_in            => s_data_in(16,6),
			data_out           => s_data_out(16,6),
			out1               => s_out1(16,6),
			out2               => s_out2(16,6),
			lock_lower_row_out => s_locks_lower_out(16,6),
			lock_lower_row_in  => s_locks_lower_in(16,6),
			in1                => s_in1(16,6),
			in2                => s_in2(16,6),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(6)
		);
	s_in1(16,6)            <= s_out1(17,6);
	s_in2(16,6)            <= s_out2(17,7);
	s_locks_lower_in(16,6) <= s_locks_lower_out(17,6);

		normal_cell_16_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,7),
			fetch              => s_fetch(16,7),
			data_in            => s_data_in(16,7),
			data_out           => s_data_out(16,7),
			out1               => s_out1(16,7),
			out2               => s_out2(16,7),
			lock_lower_row_out => s_locks_lower_out(16,7),
			lock_lower_row_in  => s_locks_lower_in(16,7),
			in1                => s_in1(16,7),
			in2                => s_in2(16,7),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(7)
		);
	s_in1(16,7)            <= s_out1(17,7);
	s_in2(16,7)            <= s_out2(17,8);
	s_locks_lower_in(16,7) <= s_locks_lower_out(17,7);

		normal_cell_16_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,8),
			fetch              => s_fetch(16,8),
			data_in            => s_data_in(16,8),
			data_out           => s_data_out(16,8),
			out1               => s_out1(16,8),
			out2               => s_out2(16,8),
			lock_lower_row_out => s_locks_lower_out(16,8),
			lock_lower_row_in  => s_locks_lower_in(16,8),
			in1                => s_in1(16,8),
			in2                => s_in2(16,8),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(8)
		);
	s_in1(16,8)            <= s_out1(17,8);
	s_in2(16,8)            <= s_out2(17,9);
	s_locks_lower_in(16,8) <= s_locks_lower_out(17,8);

		normal_cell_16_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,9),
			fetch              => s_fetch(16,9),
			data_in            => s_data_in(16,9),
			data_out           => s_data_out(16,9),
			out1               => s_out1(16,9),
			out2               => s_out2(16,9),
			lock_lower_row_out => s_locks_lower_out(16,9),
			lock_lower_row_in  => s_locks_lower_in(16,9),
			in1                => s_in1(16,9),
			in2                => s_in2(16,9),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(9)
		);
	s_in1(16,9)            <= s_out1(17,9);
	s_in2(16,9)            <= s_out2(17,10);
	s_locks_lower_in(16,9) <= s_locks_lower_out(17,9);

		normal_cell_16_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,10),
			fetch              => s_fetch(16,10),
			data_in            => s_data_in(16,10),
			data_out           => s_data_out(16,10),
			out1               => s_out1(16,10),
			out2               => s_out2(16,10),
			lock_lower_row_out => s_locks_lower_out(16,10),
			lock_lower_row_in  => s_locks_lower_in(16,10),
			in1                => s_in1(16,10),
			in2                => s_in2(16,10),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(10)
		);
	s_in1(16,10)            <= s_out1(17,10);
	s_in2(16,10)            <= s_out2(17,11);
	s_locks_lower_in(16,10) <= s_locks_lower_out(17,10);

		normal_cell_16_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,11),
			fetch              => s_fetch(16,11),
			data_in            => s_data_in(16,11),
			data_out           => s_data_out(16,11),
			out1               => s_out1(16,11),
			out2               => s_out2(16,11),
			lock_lower_row_out => s_locks_lower_out(16,11),
			lock_lower_row_in  => s_locks_lower_in(16,11),
			in1                => s_in1(16,11),
			in2                => s_in2(16,11),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(11)
		);
	s_in1(16,11)            <= s_out1(17,11);
	s_in2(16,11)            <= s_out2(17,12);
	s_locks_lower_in(16,11) <= s_locks_lower_out(17,11);

		normal_cell_16_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,12),
			fetch              => s_fetch(16,12),
			data_in            => s_data_in(16,12),
			data_out           => s_data_out(16,12),
			out1               => s_out1(16,12),
			out2               => s_out2(16,12),
			lock_lower_row_out => s_locks_lower_out(16,12),
			lock_lower_row_in  => s_locks_lower_in(16,12),
			in1                => s_in1(16,12),
			in2                => s_in2(16,12),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(12)
		);
	s_in1(16,12)            <= s_out1(17,12);
	s_in2(16,12)            <= s_out2(17,13);
	s_locks_lower_in(16,12) <= s_locks_lower_out(17,12);

		normal_cell_16_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,13),
			fetch              => s_fetch(16,13),
			data_in            => s_data_in(16,13),
			data_out           => s_data_out(16,13),
			out1               => s_out1(16,13),
			out2               => s_out2(16,13),
			lock_lower_row_out => s_locks_lower_out(16,13),
			lock_lower_row_in  => s_locks_lower_in(16,13),
			in1                => s_in1(16,13),
			in2                => s_in2(16,13),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(13)
		);
	s_in1(16,13)            <= s_out1(17,13);
	s_in2(16,13)            <= s_out2(17,14);
	s_locks_lower_in(16,13) <= s_locks_lower_out(17,13);

		normal_cell_16_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,14),
			fetch              => s_fetch(16,14),
			data_in            => s_data_in(16,14),
			data_out           => s_data_out(16,14),
			out1               => s_out1(16,14),
			out2               => s_out2(16,14),
			lock_lower_row_out => s_locks_lower_out(16,14),
			lock_lower_row_in  => s_locks_lower_in(16,14),
			in1                => s_in1(16,14),
			in2                => s_in2(16,14),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(14)
		);
	s_in1(16,14)            <= s_out1(17,14);
	s_in2(16,14)            <= s_out2(17,15);
	s_locks_lower_in(16,14) <= s_locks_lower_out(17,14);

		normal_cell_16_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,15),
			fetch              => s_fetch(16,15),
			data_in            => s_data_in(16,15),
			data_out           => s_data_out(16,15),
			out1               => s_out1(16,15),
			out2               => s_out2(16,15),
			lock_lower_row_out => s_locks_lower_out(16,15),
			lock_lower_row_in  => s_locks_lower_in(16,15),
			in1                => s_in1(16,15),
			in2                => s_in2(16,15),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(15)
		);
	s_in1(16,15)            <= s_out1(17,15);
	s_in2(16,15)            <= s_out2(17,16);
	s_locks_lower_in(16,15) <= s_locks_lower_out(17,15);

		normal_cell_16_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,16),
			fetch              => s_fetch(16,16),
			data_in            => s_data_in(16,16),
			data_out           => s_data_out(16,16),
			out1               => s_out1(16,16),
			out2               => s_out2(16,16),
			lock_lower_row_out => s_locks_lower_out(16,16),
			lock_lower_row_in  => s_locks_lower_in(16,16),
			in1                => s_in1(16,16),
			in2                => s_in2(16,16),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(16)
		);
	s_in1(16,16)            <= s_out1(17,16);
	s_in2(16,16)            <= s_out2(17,17);
	s_locks_lower_in(16,16) <= s_locks_lower_out(17,16);

		normal_cell_16_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,17),
			fetch              => s_fetch(16,17),
			data_in            => s_data_in(16,17),
			data_out           => s_data_out(16,17),
			out1               => s_out1(16,17),
			out2               => s_out2(16,17),
			lock_lower_row_out => s_locks_lower_out(16,17),
			lock_lower_row_in  => s_locks_lower_in(16,17),
			in1                => s_in1(16,17),
			in2                => s_in2(16,17),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(17)
		);
	s_in1(16,17)            <= s_out1(17,17);
	s_in2(16,17)            <= s_out2(17,18);
	s_locks_lower_in(16,17) <= s_locks_lower_out(17,17);

		normal_cell_16_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,18),
			fetch              => s_fetch(16,18),
			data_in            => s_data_in(16,18),
			data_out           => s_data_out(16,18),
			out1               => s_out1(16,18),
			out2               => s_out2(16,18),
			lock_lower_row_out => s_locks_lower_out(16,18),
			lock_lower_row_in  => s_locks_lower_in(16,18),
			in1                => s_in1(16,18),
			in2                => s_in2(16,18),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(18)
		);
	s_in1(16,18)            <= s_out1(17,18);
	s_in2(16,18)            <= s_out2(17,19);
	s_locks_lower_in(16,18) <= s_locks_lower_out(17,18);

		normal_cell_16_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,19),
			fetch              => s_fetch(16,19),
			data_in            => s_data_in(16,19),
			data_out           => s_data_out(16,19),
			out1               => s_out1(16,19),
			out2               => s_out2(16,19),
			lock_lower_row_out => s_locks_lower_out(16,19),
			lock_lower_row_in  => s_locks_lower_in(16,19),
			in1                => s_in1(16,19),
			in2                => s_in2(16,19),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(19)
		);
	s_in1(16,19)            <= s_out1(17,19);
	s_in2(16,19)            <= s_out2(17,20);
	s_locks_lower_in(16,19) <= s_locks_lower_out(17,19);

		normal_cell_16_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,20),
			fetch              => s_fetch(16,20),
			data_in            => s_data_in(16,20),
			data_out           => s_data_out(16,20),
			out1               => s_out1(16,20),
			out2               => s_out2(16,20),
			lock_lower_row_out => s_locks_lower_out(16,20),
			lock_lower_row_in  => s_locks_lower_in(16,20),
			in1                => s_in1(16,20),
			in2                => s_in2(16,20),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(20)
		);
	s_in1(16,20)            <= s_out1(17,20);
	s_in2(16,20)            <= s_out2(17,21);
	s_locks_lower_in(16,20) <= s_locks_lower_out(17,20);

		normal_cell_16_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,21),
			fetch              => s_fetch(16,21),
			data_in            => s_data_in(16,21),
			data_out           => s_data_out(16,21),
			out1               => s_out1(16,21),
			out2               => s_out2(16,21),
			lock_lower_row_out => s_locks_lower_out(16,21),
			lock_lower_row_in  => s_locks_lower_in(16,21),
			in1                => s_in1(16,21),
			in2                => s_in2(16,21),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(21)
		);
	s_in1(16,21)            <= s_out1(17,21);
	s_in2(16,21)            <= s_out2(17,22);
	s_locks_lower_in(16,21) <= s_locks_lower_out(17,21);

		normal_cell_16_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,22),
			fetch              => s_fetch(16,22),
			data_in            => s_data_in(16,22),
			data_out           => s_data_out(16,22),
			out1               => s_out1(16,22),
			out2               => s_out2(16,22),
			lock_lower_row_out => s_locks_lower_out(16,22),
			lock_lower_row_in  => s_locks_lower_in(16,22),
			in1                => s_in1(16,22),
			in2                => s_in2(16,22),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(22)
		);
	s_in1(16,22)            <= s_out1(17,22);
	s_in2(16,22)            <= s_out2(17,23);
	s_locks_lower_in(16,22) <= s_locks_lower_out(17,22);

		normal_cell_16_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,23),
			fetch              => s_fetch(16,23),
			data_in            => s_data_in(16,23),
			data_out           => s_data_out(16,23),
			out1               => s_out1(16,23),
			out2               => s_out2(16,23),
			lock_lower_row_out => s_locks_lower_out(16,23),
			lock_lower_row_in  => s_locks_lower_in(16,23),
			in1                => s_in1(16,23),
			in2                => s_in2(16,23),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(23)
		);
	s_in1(16,23)            <= s_out1(17,23);
	s_in2(16,23)            <= s_out2(17,24);
	s_locks_lower_in(16,23) <= s_locks_lower_out(17,23);

		normal_cell_16_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,24),
			fetch              => s_fetch(16,24),
			data_in            => s_data_in(16,24),
			data_out           => s_data_out(16,24),
			out1               => s_out1(16,24),
			out2               => s_out2(16,24),
			lock_lower_row_out => s_locks_lower_out(16,24),
			lock_lower_row_in  => s_locks_lower_in(16,24),
			in1                => s_in1(16,24),
			in2                => s_in2(16,24),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(24)
		);
	s_in1(16,24)            <= s_out1(17,24);
	s_in2(16,24)            <= s_out2(17,25);
	s_locks_lower_in(16,24) <= s_locks_lower_out(17,24);

		normal_cell_16_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,25),
			fetch              => s_fetch(16,25),
			data_in            => s_data_in(16,25),
			data_out           => s_data_out(16,25),
			out1               => s_out1(16,25),
			out2               => s_out2(16,25),
			lock_lower_row_out => s_locks_lower_out(16,25),
			lock_lower_row_in  => s_locks_lower_in(16,25),
			in1                => s_in1(16,25),
			in2                => s_in2(16,25),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(25)
		);
	s_in1(16,25)            <= s_out1(17,25);
	s_in2(16,25)            <= s_out2(17,26);
	s_locks_lower_in(16,25) <= s_locks_lower_out(17,25);

		normal_cell_16_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,26),
			fetch              => s_fetch(16,26),
			data_in            => s_data_in(16,26),
			data_out           => s_data_out(16,26),
			out1               => s_out1(16,26),
			out2               => s_out2(16,26),
			lock_lower_row_out => s_locks_lower_out(16,26),
			lock_lower_row_in  => s_locks_lower_in(16,26),
			in1                => s_in1(16,26),
			in2                => s_in2(16,26),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(26)
		);
	s_in1(16,26)            <= s_out1(17,26);
	s_in2(16,26)            <= s_out2(17,27);
	s_locks_lower_in(16,26) <= s_locks_lower_out(17,26);

		normal_cell_16_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,27),
			fetch              => s_fetch(16,27),
			data_in            => s_data_in(16,27),
			data_out           => s_data_out(16,27),
			out1               => s_out1(16,27),
			out2               => s_out2(16,27),
			lock_lower_row_out => s_locks_lower_out(16,27),
			lock_lower_row_in  => s_locks_lower_in(16,27),
			in1                => s_in1(16,27),
			in2                => s_in2(16,27),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(27)
		);
	s_in1(16,27)            <= s_out1(17,27);
	s_in2(16,27)            <= s_out2(17,28);
	s_locks_lower_in(16,27) <= s_locks_lower_out(17,27);

		normal_cell_16_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,28),
			fetch              => s_fetch(16,28),
			data_in            => s_data_in(16,28),
			data_out           => s_data_out(16,28),
			out1               => s_out1(16,28),
			out2               => s_out2(16,28),
			lock_lower_row_out => s_locks_lower_out(16,28),
			lock_lower_row_in  => s_locks_lower_in(16,28),
			in1                => s_in1(16,28),
			in2                => s_in2(16,28),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(28)
		);
	s_in1(16,28)            <= s_out1(17,28);
	s_in2(16,28)            <= s_out2(17,29);
	s_locks_lower_in(16,28) <= s_locks_lower_out(17,28);

		normal_cell_16_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,29),
			fetch              => s_fetch(16,29),
			data_in            => s_data_in(16,29),
			data_out           => s_data_out(16,29),
			out1               => s_out1(16,29),
			out2               => s_out2(16,29),
			lock_lower_row_out => s_locks_lower_out(16,29),
			lock_lower_row_in  => s_locks_lower_in(16,29),
			in1                => s_in1(16,29),
			in2                => s_in2(16,29),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(29)
		);
	s_in1(16,29)            <= s_out1(17,29);
	s_in2(16,29)            <= s_out2(17,30);
	s_locks_lower_in(16,29) <= s_locks_lower_out(17,29);

		normal_cell_16_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,30),
			fetch              => s_fetch(16,30),
			data_in            => s_data_in(16,30),
			data_out           => s_data_out(16,30),
			out1               => s_out1(16,30),
			out2               => s_out2(16,30),
			lock_lower_row_out => s_locks_lower_out(16,30),
			lock_lower_row_in  => s_locks_lower_in(16,30),
			in1                => s_in1(16,30),
			in2                => s_in2(16,30),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(30)
		);
	s_in1(16,30)            <= s_out1(17,30);
	s_in2(16,30)            <= s_out2(17,31);
	s_locks_lower_in(16,30) <= s_locks_lower_out(17,30);

		normal_cell_16_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,31),
			fetch              => s_fetch(16,31),
			data_in            => s_data_in(16,31),
			data_out           => s_data_out(16,31),
			out1               => s_out1(16,31),
			out2               => s_out2(16,31),
			lock_lower_row_out => s_locks_lower_out(16,31),
			lock_lower_row_in  => s_locks_lower_in(16,31),
			in1                => s_in1(16,31),
			in2                => s_in2(16,31),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(31)
		);
	s_in1(16,31)            <= s_out1(17,31);
	s_in2(16,31)            <= s_out2(17,32);
	s_locks_lower_in(16,31) <= s_locks_lower_out(17,31);

		normal_cell_16_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,32),
			fetch              => s_fetch(16,32),
			data_in            => s_data_in(16,32),
			data_out           => s_data_out(16,32),
			out1               => s_out1(16,32),
			out2               => s_out2(16,32),
			lock_lower_row_out => s_locks_lower_out(16,32),
			lock_lower_row_in  => s_locks_lower_in(16,32),
			in1                => s_in1(16,32),
			in2                => s_in2(16,32),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(32)
		);
	s_in1(16,32)            <= s_out1(17,32);
	s_in2(16,32)            <= s_out2(17,33);
	s_locks_lower_in(16,32) <= s_locks_lower_out(17,32);

		normal_cell_16_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,33),
			fetch              => s_fetch(16,33),
			data_in            => s_data_in(16,33),
			data_out           => s_data_out(16,33),
			out1               => s_out1(16,33),
			out2               => s_out2(16,33),
			lock_lower_row_out => s_locks_lower_out(16,33),
			lock_lower_row_in  => s_locks_lower_in(16,33),
			in1                => s_in1(16,33),
			in2                => s_in2(16,33),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(33)
		);
	s_in1(16,33)            <= s_out1(17,33);
	s_in2(16,33)            <= s_out2(17,34);
	s_locks_lower_in(16,33) <= s_locks_lower_out(17,33);

		normal_cell_16_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,34),
			fetch              => s_fetch(16,34),
			data_in            => s_data_in(16,34),
			data_out           => s_data_out(16,34),
			out1               => s_out1(16,34),
			out2               => s_out2(16,34),
			lock_lower_row_out => s_locks_lower_out(16,34),
			lock_lower_row_in  => s_locks_lower_in(16,34),
			in1                => s_in1(16,34),
			in2                => s_in2(16,34),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(34)
		);
	s_in1(16,34)            <= s_out1(17,34);
	s_in2(16,34)            <= s_out2(17,35);
	s_locks_lower_in(16,34) <= s_locks_lower_out(17,34);

		normal_cell_16_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,35),
			fetch              => s_fetch(16,35),
			data_in            => s_data_in(16,35),
			data_out           => s_data_out(16,35),
			out1               => s_out1(16,35),
			out2               => s_out2(16,35),
			lock_lower_row_out => s_locks_lower_out(16,35),
			lock_lower_row_in  => s_locks_lower_in(16,35),
			in1                => s_in1(16,35),
			in2                => s_in2(16,35),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(35)
		);
	s_in1(16,35)            <= s_out1(17,35);
	s_in2(16,35)            <= s_out2(17,36);
	s_locks_lower_in(16,35) <= s_locks_lower_out(17,35);

		normal_cell_16_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,36),
			fetch              => s_fetch(16,36),
			data_in            => s_data_in(16,36),
			data_out           => s_data_out(16,36),
			out1               => s_out1(16,36),
			out2               => s_out2(16,36),
			lock_lower_row_out => s_locks_lower_out(16,36),
			lock_lower_row_in  => s_locks_lower_in(16,36),
			in1                => s_in1(16,36),
			in2                => s_in2(16,36),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(36)
		);
	s_in1(16,36)            <= s_out1(17,36);
	s_in2(16,36)            <= s_out2(17,37);
	s_locks_lower_in(16,36) <= s_locks_lower_out(17,36);

		normal_cell_16_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,37),
			fetch              => s_fetch(16,37),
			data_in            => s_data_in(16,37),
			data_out           => s_data_out(16,37),
			out1               => s_out1(16,37),
			out2               => s_out2(16,37),
			lock_lower_row_out => s_locks_lower_out(16,37),
			lock_lower_row_in  => s_locks_lower_in(16,37),
			in1                => s_in1(16,37),
			in2                => s_in2(16,37),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(37)
		);
	s_in1(16,37)            <= s_out1(17,37);
	s_in2(16,37)            <= s_out2(17,38);
	s_locks_lower_in(16,37) <= s_locks_lower_out(17,37);

		normal_cell_16_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,38),
			fetch              => s_fetch(16,38),
			data_in            => s_data_in(16,38),
			data_out           => s_data_out(16,38),
			out1               => s_out1(16,38),
			out2               => s_out2(16,38),
			lock_lower_row_out => s_locks_lower_out(16,38),
			lock_lower_row_in  => s_locks_lower_in(16,38),
			in1                => s_in1(16,38),
			in2                => s_in2(16,38),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(38)
		);
	s_in1(16,38)            <= s_out1(17,38);
	s_in2(16,38)            <= s_out2(17,39);
	s_locks_lower_in(16,38) <= s_locks_lower_out(17,38);

		normal_cell_16_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,39),
			fetch              => s_fetch(16,39),
			data_in            => s_data_in(16,39),
			data_out           => s_data_out(16,39),
			out1               => s_out1(16,39),
			out2               => s_out2(16,39),
			lock_lower_row_out => s_locks_lower_out(16,39),
			lock_lower_row_in  => s_locks_lower_in(16,39),
			in1                => s_in1(16,39),
			in2                => s_in2(16,39),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(39)
		);
	s_in1(16,39)            <= s_out1(17,39);
	s_in2(16,39)            <= s_out2(17,40);
	s_locks_lower_in(16,39) <= s_locks_lower_out(17,39);

		normal_cell_16_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,40),
			fetch              => s_fetch(16,40),
			data_in            => s_data_in(16,40),
			data_out           => s_data_out(16,40),
			out1               => s_out1(16,40),
			out2               => s_out2(16,40),
			lock_lower_row_out => s_locks_lower_out(16,40),
			lock_lower_row_in  => s_locks_lower_in(16,40),
			in1                => s_in1(16,40),
			in2                => s_in2(16,40),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(40)
		);
	s_in1(16,40)            <= s_out1(17,40);
	s_in2(16,40)            <= s_out2(17,41);
	s_locks_lower_in(16,40) <= s_locks_lower_out(17,40);

		normal_cell_16_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,41),
			fetch              => s_fetch(16,41),
			data_in            => s_data_in(16,41),
			data_out           => s_data_out(16,41),
			out1               => s_out1(16,41),
			out2               => s_out2(16,41),
			lock_lower_row_out => s_locks_lower_out(16,41),
			lock_lower_row_in  => s_locks_lower_in(16,41),
			in1                => s_in1(16,41),
			in2                => s_in2(16,41),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(41)
		);
	s_in1(16,41)            <= s_out1(17,41);
	s_in2(16,41)            <= s_out2(17,42);
	s_locks_lower_in(16,41) <= s_locks_lower_out(17,41);

		normal_cell_16_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,42),
			fetch              => s_fetch(16,42),
			data_in            => s_data_in(16,42),
			data_out           => s_data_out(16,42),
			out1               => s_out1(16,42),
			out2               => s_out2(16,42),
			lock_lower_row_out => s_locks_lower_out(16,42),
			lock_lower_row_in  => s_locks_lower_in(16,42),
			in1                => s_in1(16,42),
			in2                => s_in2(16,42),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(42)
		);
	s_in1(16,42)            <= s_out1(17,42);
	s_in2(16,42)            <= s_out2(17,43);
	s_locks_lower_in(16,42) <= s_locks_lower_out(17,42);

		normal_cell_16_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,43),
			fetch              => s_fetch(16,43),
			data_in            => s_data_in(16,43),
			data_out           => s_data_out(16,43),
			out1               => s_out1(16,43),
			out2               => s_out2(16,43),
			lock_lower_row_out => s_locks_lower_out(16,43),
			lock_lower_row_in  => s_locks_lower_in(16,43),
			in1                => s_in1(16,43),
			in2                => s_in2(16,43),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(43)
		);
	s_in1(16,43)            <= s_out1(17,43);
	s_in2(16,43)            <= s_out2(17,44);
	s_locks_lower_in(16,43) <= s_locks_lower_out(17,43);

		normal_cell_16_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,44),
			fetch              => s_fetch(16,44),
			data_in            => s_data_in(16,44),
			data_out           => s_data_out(16,44),
			out1               => s_out1(16,44),
			out2               => s_out2(16,44),
			lock_lower_row_out => s_locks_lower_out(16,44),
			lock_lower_row_in  => s_locks_lower_in(16,44),
			in1                => s_in1(16,44),
			in2                => s_in2(16,44),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(44)
		);
	s_in1(16,44)            <= s_out1(17,44);
	s_in2(16,44)            <= s_out2(17,45);
	s_locks_lower_in(16,44) <= s_locks_lower_out(17,44);

		normal_cell_16_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,45),
			fetch              => s_fetch(16,45),
			data_in            => s_data_in(16,45),
			data_out           => s_data_out(16,45),
			out1               => s_out1(16,45),
			out2               => s_out2(16,45),
			lock_lower_row_out => s_locks_lower_out(16,45),
			lock_lower_row_in  => s_locks_lower_in(16,45),
			in1                => s_in1(16,45),
			in2                => s_in2(16,45),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(45)
		);
	s_in1(16,45)            <= s_out1(17,45);
	s_in2(16,45)            <= s_out2(17,46);
	s_locks_lower_in(16,45) <= s_locks_lower_out(17,45);

		normal_cell_16_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,46),
			fetch              => s_fetch(16,46),
			data_in            => s_data_in(16,46),
			data_out           => s_data_out(16,46),
			out1               => s_out1(16,46),
			out2               => s_out2(16,46),
			lock_lower_row_out => s_locks_lower_out(16,46),
			lock_lower_row_in  => s_locks_lower_in(16,46),
			in1                => s_in1(16,46),
			in2                => s_in2(16,46),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(46)
		);
	s_in1(16,46)            <= s_out1(17,46);
	s_in2(16,46)            <= s_out2(17,47);
	s_locks_lower_in(16,46) <= s_locks_lower_out(17,46);

		normal_cell_16_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,47),
			fetch              => s_fetch(16,47),
			data_in            => s_data_in(16,47),
			data_out           => s_data_out(16,47),
			out1               => s_out1(16,47),
			out2               => s_out2(16,47),
			lock_lower_row_out => s_locks_lower_out(16,47),
			lock_lower_row_in  => s_locks_lower_in(16,47),
			in1                => s_in1(16,47),
			in2                => s_in2(16,47),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(47)
		);
	s_in1(16,47)            <= s_out1(17,47);
	s_in2(16,47)            <= s_out2(17,48);
	s_locks_lower_in(16,47) <= s_locks_lower_out(17,47);

		normal_cell_16_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,48),
			fetch              => s_fetch(16,48),
			data_in            => s_data_in(16,48),
			data_out           => s_data_out(16,48),
			out1               => s_out1(16,48),
			out2               => s_out2(16,48),
			lock_lower_row_out => s_locks_lower_out(16,48),
			lock_lower_row_in  => s_locks_lower_in(16,48),
			in1                => s_in1(16,48),
			in2                => s_in2(16,48),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(48)
		);
	s_in1(16,48)            <= s_out1(17,48);
	s_in2(16,48)            <= s_out2(17,49);
	s_locks_lower_in(16,48) <= s_locks_lower_out(17,48);

		normal_cell_16_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,49),
			fetch              => s_fetch(16,49),
			data_in            => s_data_in(16,49),
			data_out           => s_data_out(16,49),
			out1               => s_out1(16,49),
			out2               => s_out2(16,49),
			lock_lower_row_out => s_locks_lower_out(16,49),
			lock_lower_row_in  => s_locks_lower_in(16,49),
			in1                => s_in1(16,49),
			in2                => s_in2(16,49),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(49)
		);
	s_in1(16,49)            <= s_out1(17,49);
	s_in2(16,49)            <= s_out2(17,50);
	s_locks_lower_in(16,49) <= s_locks_lower_out(17,49);

		normal_cell_16_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,50),
			fetch              => s_fetch(16,50),
			data_in            => s_data_in(16,50),
			data_out           => s_data_out(16,50),
			out1               => s_out1(16,50),
			out2               => s_out2(16,50),
			lock_lower_row_out => s_locks_lower_out(16,50),
			lock_lower_row_in  => s_locks_lower_in(16,50),
			in1                => s_in1(16,50),
			in2                => s_in2(16,50),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(50)
		);
	s_in1(16,50)            <= s_out1(17,50);
	s_in2(16,50)            <= s_out2(17,51);
	s_locks_lower_in(16,50) <= s_locks_lower_out(17,50);

		normal_cell_16_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,51),
			fetch              => s_fetch(16,51),
			data_in            => s_data_in(16,51),
			data_out           => s_data_out(16,51),
			out1               => s_out1(16,51),
			out2               => s_out2(16,51),
			lock_lower_row_out => s_locks_lower_out(16,51),
			lock_lower_row_in  => s_locks_lower_in(16,51),
			in1                => s_in1(16,51),
			in2                => s_in2(16,51),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(51)
		);
	s_in1(16,51)            <= s_out1(17,51);
	s_in2(16,51)            <= s_out2(17,52);
	s_locks_lower_in(16,51) <= s_locks_lower_out(17,51);

		normal_cell_16_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,52),
			fetch              => s_fetch(16,52),
			data_in            => s_data_in(16,52),
			data_out           => s_data_out(16,52),
			out1               => s_out1(16,52),
			out2               => s_out2(16,52),
			lock_lower_row_out => s_locks_lower_out(16,52),
			lock_lower_row_in  => s_locks_lower_in(16,52),
			in1                => s_in1(16,52),
			in2                => s_in2(16,52),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(52)
		);
	s_in1(16,52)            <= s_out1(17,52);
	s_in2(16,52)            <= s_out2(17,53);
	s_locks_lower_in(16,52) <= s_locks_lower_out(17,52);

		normal_cell_16_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,53),
			fetch              => s_fetch(16,53),
			data_in            => s_data_in(16,53),
			data_out           => s_data_out(16,53),
			out1               => s_out1(16,53),
			out2               => s_out2(16,53),
			lock_lower_row_out => s_locks_lower_out(16,53),
			lock_lower_row_in  => s_locks_lower_in(16,53),
			in1                => s_in1(16,53),
			in2                => s_in2(16,53),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(53)
		);
	s_in1(16,53)            <= s_out1(17,53);
	s_in2(16,53)            <= s_out2(17,54);
	s_locks_lower_in(16,53) <= s_locks_lower_out(17,53);

		normal_cell_16_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,54),
			fetch              => s_fetch(16,54),
			data_in            => s_data_in(16,54),
			data_out           => s_data_out(16,54),
			out1               => s_out1(16,54),
			out2               => s_out2(16,54),
			lock_lower_row_out => s_locks_lower_out(16,54),
			lock_lower_row_in  => s_locks_lower_in(16,54),
			in1                => s_in1(16,54),
			in2                => s_in2(16,54),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(54)
		);
	s_in1(16,54)            <= s_out1(17,54);
	s_in2(16,54)            <= s_out2(17,55);
	s_locks_lower_in(16,54) <= s_locks_lower_out(17,54);

		normal_cell_16_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,55),
			fetch              => s_fetch(16,55),
			data_in            => s_data_in(16,55),
			data_out           => s_data_out(16,55),
			out1               => s_out1(16,55),
			out2               => s_out2(16,55),
			lock_lower_row_out => s_locks_lower_out(16,55),
			lock_lower_row_in  => s_locks_lower_in(16,55),
			in1                => s_in1(16,55),
			in2                => s_in2(16,55),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(55)
		);
	s_in1(16,55)            <= s_out1(17,55);
	s_in2(16,55)            <= s_out2(17,56);
	s_locks_lower_in(16,55) <= s_locks_lower_out(17,55);

		normal_cell_16_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,56),
			fetch              => s_fetch(16,56),
			data_in            => s_data_in(16,56),
			data_out           => s_data_out(16,56),
			out1               => s_out1(16,56),
			out2               => s_out2(16,56),
			lock_lower_row_out => s_locks_lower_out(16,56),
			lock_lower_row_in  => s_locks_lower_in(16,56),
			in1                => s_in1(16,56),
			in2                => s_in2(16,56),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(56)
		);
	s_in1(16,56)            <= s_out1(17,56);
	s_in2(16,56)            <= s_out2(17,57);
	s_locks_lower_in(16,56) <= s_locks_lower_out(17,56);

		normal_cell_16_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,57),
			fetch              => s_fetch(16,57),
			data_in            => s_data_in(16,57),
			data_out           => s_data_out(16,57),
			out1               => s_out1(16,57),
			out2               => s_out2(16,57),
			lock_lower_row_out => s_locks_lower_out(16,57),
			lock_lower_row_in  => s_locks_lower_in(16,57),
			in1                => s_in1(16,57),
			in2                => s_in2(16,57),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(57)
		);
	s_in1(16,57)            <= s_out1(17,57);
	s_in2(16,57)            <= s_out2(17,58);
	s_locks_lower_in(16,57) <= s_locks_lower_out(17,57);

		normal_cell_16_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,58),
			fetch              => s_fetch(16,58),
			data_in            => s_data_in(16,58),
			data_out           => s_data_out(16,58),
			out1               => s_out1(16,58),
			out2               => s_out2(16,58),
			lock_lower_row_out => s_locks_lower_out(16,58),
			lock_lower_row_in  => s_locks_lower_in(16,58),
			in1                => s_in1(16,58),
			in2                => s_in2(16,58),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(58)
		);
	s_in1(16,58)            <= s_out1(17,58);
	s_in2(16,58)            <= s_out2(17,59);
	s_locks_lower_in(16,58) <= s_locks_lower_out(17,58);

		normal_cell_16_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,59),
			fetch              => s_fetch(16,59),
			data_in            => s_data_in(16,59),
			data_out           => s_data_out(16,59),
			out1               => s_out1(16,59),
			out2               => s_out2(16,59),
			lock_lower_row_out => s_locks_lower_out(16,59),
			lock_lower_row_in  => s_locks_lower_in(16,59),
			in1                => s_in1(16,59),
			in2                => s_in2(16,59),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(59)
		);
	s_in1(16,59)            <= s_out1(17,59);
	s_in2(16,59)            <= s_out2(17,60);
	s_locks_lower_in(16,59) <= s_locks_lower_out(17,59);

		last_col_cell_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(16,60),
			fetch              => s_fetch(16,60),
			data_in            => s_data_in(16,60),
			data_out           => s_data_out(16,60),
			out1               => s_out1(16,60),
			out2               => s_out2(16,60),
			lock_lower_row_out => s_locks_lower_out(16,60),
			lock_lower_row_in  => s_locks_lower_in(16,60),
			in1                => s_in1(16,60),
			in2                => (others => '0'),
			lock_row           => s_locks(16),
			piv_found          => s_piv_found,
			row_data           => s_row_data(16),
			col_data           => s_col_data(60)
		);
	s_in1(16,60)            <= s_out1(17,60);
	s_locks_lower_in(16,60) <= s_locks_lower_out(17,60);

		normal_cell_17_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,1),
			fetch              => s_fetch(17,1),
			data_in            => s_data_in(17,1),
			data_out           => s_data_out(17,1),
			out1               => s_out1(17,1),
			out2               => s_out2(17,1),
			lock_lower_row_out => s_locks_lower_out(17,1),
			lock_lower_row_in  => s_locks_lower_in(17,1),
			in1                => s_in1(17,1),
			in2                => s_in2(17,1),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(1)
		);
	s_in1(17,1)            <= s_out1(18,1);
	s_in2(17,1)            <= s_out2(18,2);
	s_locks_lower_in(17,1) <= s_locks_lower_out(18,1);

		normal_cell_17_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,2),
			fetch              => s_fetch(17,2),
			data_in            => s_data_in(17,2),
			data_out           => s_data_out(17,2),
			out1               => s_out1(17,2),
			out2               => s_out2(17,2),
			lock_lower_row_out => s_locks_lower_out(17,2),
			lock_lower_row_in  => s_locks_lower_in(17,2),
			in1                => s_in1(17,2),
			in2                => s_in2(17,2),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(2)
		);
	s_in1(17,2)            <= s_out1(18,2);
	s_in2(17,2)            <= s_out2(18,3);
	s_locks_lower_in(17,2) <= s_locks_lower_out(18,2);

		normal_cell_17_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,3),
			fetch              => s_fetch(17,3),
			data_in            => s_data_in(17,3),
			data_out           => s_data_out(17,3),
			out1               => s_out1(17,3),
			out2               => s_out2(17,3),
			lock_lower_row_out => s_locks_lower_out(17,3),
			lock_lower_row_in  => s_locks_lower_in(17,3),
			in1                => s_in1(17,3),
			in2                => s_in2(17,3),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(3)
		);
	s_in1(17,3)            <= s_out1(18,3);
	s_in2(17,3)            <= s_out2(18,4);
	s_locks_lower_in(17,3) <= s_locks_lower_out(18,3);

		normal_cell_17_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,4),
			fetch              => s_fetch(17,4),
			data_in            => s_data_in(17,4),
			data_out           => s_data_out(17,4),
			out1               => s_out1(17,4),
			out2               => s_out2(17,4),
			lock_lower_row_out => s_locks_lower_out(17,4),
			lock_lower_row_in  => s_locks_lower_in(17,4),
			in1                => s_in1(17,4),
			in2                => s_in2(17,4),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(4)
		);
	s_in1(17,4)            <= s_out1(18,4);
	s_in2(17,4)            <= s_out2(18,5);
	s_locks_lower_in(17,4) <= s_locks_lower_out(18,4);

		normal_cell_17_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,5),
			fetch              => s_fetch(17,5),
			data_in            => s_data_in(17,5),
			data_out           => s_data_out(17,5),
			out1               => s_out1(17,5),
			out2               => s_out2(17,5),
			lock_lower_row_out => s_locks_lower_out(17,5),
			lock_lower_row_in  => s_locks_lower_in(17,5),
			in1                => s_in1(17,5),
			in2                => s_in2(17,5),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(5)
		);
	s_in1(17,5)            <= s_out1(18,5);
	s_in2(17,5)            <= s_out2(18,6);
	s_locks_lower_in(17,5) <= s_locks_lower_out(18,5);

		normal_cell_17_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,6),
			fetch              => s_fetch(17,6),
			data_in            => s_data_in(17,6),
			data_out           => s_data_out(17,6),
			out1               => s_out1(17,6),
			out2               => s_out2(17,6),
			lock_lower_row_out => s_locks_lower_out(17,6),
			lock_lower_row_in  => s_locks_lower_in(17,6),
			in1                => s_in1(17,6),
			in2                => s_in2(17,6),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(6)
		);
	s_in1(17,6)            <= s_out1(18,6);
	s_in2(17,6)            <= s_out2(18,7);
	s_locks_lower_in(17,6) <= s_locks_lower_out(18,6);

		normal_cell_17_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,7),
			fetch              => s_fetch(17,7),
			data_in            => s_data_in(17,7),
			data_out           => s_data_out(17,7),
			out1               => s_out1(17,7),
			out2               => s_out2(17,7),
			lock_lower_row_out => s_locks_lower_out(17,7),
			lock_lower_row_in  => s_locks_lower_in(17,7),
			in1                => s_in1(17,7),
			in2                => s_in2(17,7),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(7)
		);
	s_in1(17,7)            <= s_out1(18,7);
	s_in2(17,7)            <= s_out2(18,8);
	s_locks_lower_in(17,7) <= s_locks_lower_out(18,7);

		normal_cell_17_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,8),
			fetch              => s_fetch(17,8),
			data_in            => s_data_in(17,8),
			data_out           => s_data_out(17,8),
			out1               => s_out1(17,8),
			out2               => s_out2(17,8),
			lock_lower_row_out => s_locks_lower_out(17,8),
			lock_lower_row_in  => s_locks_lower_in(17,8),
			in1                => s_in1(17,8),
			in2                => s_in2(17,8),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(8)
		);
	s_in1(17,8)            <= s_out1(18,8);
	s_in2(17,8)            <= s_out2(18,9);
	s_locks_lower_in(17,8) <= s_locks_lower_out(18,8);

		normal_cell_17_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,9),
			fetch              => s_fetch(17,9),
			data_in            => s_data_in(17,9),
			data_out           => s_data_out(17,9),
			out1               => s_out1(17,9),
			out2               => s_out2(17,9),
			lock_lower_row_out => s_locks_lower_out(17,9),
			lock_lower_row_in  => s_locks_lower_in(17,9),
			in1                => s_in1(17,9),
			in2                => s_in2(17,9),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(9)
		);
	s_in1(17,9)            <= s_out1(18,9);
	s_in2(17,9)            <= s_out2(18,10);
	s_locks_lower_in(17,9) <= s_locks_lower_out(18,9);

		normal_cell_17_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,10),
			fetch              => s_fetch(17,10),
			data_in            => s_data_in(17,10),
			data_out           => s_data_out(17,10),
			out1               => s_out1(17,10),
			out2               => s_out2(17,10),
			lock_lower_row_out => s_locks_lower_out(17,10),
			lock_lower_row_in  => s_locks_lower_in(17,10),
			in1                => s_in1(17,10),
			in2                => s_in2(17,10),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(10)
		);
	s_in1(17,10)            <= s_out1(18,10);
	s_in2(17,10)            <= s_out2(18,11);
	s_locks_lower_in(17,10) <= s_locks_lower_out(18,10);

		normal_cell_17_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,11),
			fetch              => s_fetch(17,11),
			data_in            => s_data_in(17,11),
			data_out           => s_data_out(17,11),
			out1               => s_out1(17,11),
			out2               => s_out2(17,11),
			lock_lower_row_out => s_locks_lower_out(17,11),
			lock_lower_row_in  => s_locks_lower_in(17,11),
			in1                => s_in1(17,11),
			in2                => s_in2(17,11),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(11)
		);
	s_in1(17,11)            <= s_out1(18,11);
	s_in2(17,11)            <= s_out2(18,12);
	s_locks_lower_in(17,11) <= s_locks_lower_out(18,11);

		normal_cell_17_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,12),
			fetch              => s_fetch(17,12),
			data_in            => s_data_in(17,12),
			data_out           => s_data_out(17,12),
			out1               => s_out1(17,12),
			out2               => s_out2(17,12),
			lock_lower_row_out => s_locks_lower_out(17,12),
			lock_lower_row_in  => s_locks_lower_in(17,12),
			in1                => s_in1(17,12),
			in2                => s_in2(17,12),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(12)
		);
	s_in1(17,12)            <= s_out1(18,12);
	s_in2(17,12)            <= s_out2(18,13);
	s_locks_lower_in(17,12) <= s_locks_lower_out(18,12);

		normal_cell_17_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,13),
			fetch              => s_fetch(17,13),
			data_in            => s_data_in(17,13),
			data_out           => s_data_out(17,13),
			out1               => s_out1(17,13),
			out2               => s_out2(17,13),
			lock_lower_row_out => s_locks_lower_out(17,13),
			lock_lower_row_in  => s_locks_lower_in(17,13),
			in1                => s_in1(17,13),
			in2                => s_in2(17,13),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(13)
		);
	s_in1(17,13)            <= s_out1(18,13);
	s_in2(17,13)            <= s_out2(18,14);
	s_locks_lower_in(17,13) <= s_locks_lower_out(18,13);

		normal_cell_17_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,14),
			fetch              => s_fetch(17,14),
			data_in            => s_data_in(17,14),
			data_out           => s_data_out(17,14),
			out1               => s_out1(17,14),
			out2               => s_out2(17,14),
			lock_lower_row_out => s_locks_lower_out(17,14),
			lock_lower_row_in  => s_locks_lower_in(17,14),
			in1                => s_in1(17,14),
			in2                => s_in2(17,14),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(14)
		);
	s_in1(17,14)            <= s_out1(18,14);
	s_in2(17,14)            <= s_out2(18,15);
	s_locks_lower_in(17,14) <= s_locks_lower_out(18,14);

		normal_cell_17_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,15),
			fetch              => s_fetch(17,15),
			data_in            => s_data_in(17,15),
			data_out           => s_data_out(17,15),
			out1               => s_out1(17,15),
			out2               => s_out2(17,15),
			lock_lower_row_out => s_locks_lower_out(17,15),
			lock_lower_row_in  => s_locks_lower_in(17,15),
			in1                => s_in1(17,15),
			in2                => s_in2(17,15),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(15)
		);
	s_in1(17,15)            <= s_out1(18,15);
	s_in2(17,15)            <= s_out2(18,16);
	s_locks_lower_in(17,15) <= s_locks_lower_out(18,15);

		normal_cell_17_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,16),
			fetch              => s_fetch(17,16),
			data_in            => s_data_in(17,16),
			data_out           => s_data_out(17,16),
			out1               => s_out1(17,16),
			out2               => s_out2(17,16),
			lock_lower_row_out => s_locks_lower_out(17,16),
			lock_lower_row_in  => s_locks_lower_in(17,16),
			in1                => s_in1(17,16),
			in2                => s_in2(17,16),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(16)
		);
	s_in1(17,16)            <= s_out1(18,16);
	s_in2(17,16)            <= s_out2(18,17);
	s_locks_lower_in(17,16) <= s_locks_lower_out(18,16);

		normal_cell_17_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,17),
			fetch              => s_fetch(17,17),
			data_in            => s_data_in(17,17),
			data_out           => s_data_out(17,17),
			out1               => s_out1(17,17),
			out2               => s_out2(17,17),
			lock_lower_row_out => s_locks_lower_out(17,17),
			lock_lower_row_in  => s_locks_lower_in(17,17),
			in1                => s_in1(17,17),
			in2                => s_in2(17,17),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(17)
		);
	s_in1(17,17)            <= s_out1(18,17);
	s_in2(17,17)            <= s_out2(18,18);
	s_locks_lower_in(17,17) <= s_locks_lower_out(18,17);

		normal_cell_17_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,18),
			fetch              => s_fetch(17,18),
			data_in            => s_data_in(17,18),
			data_out           => s_data_out(17,18),
			out1               => s_out1(17,18),
			out2               => s_out2(17,18),
			lock_lower_row_out => s_locks_lower_out(17,18),
			lock_lower_row_in  => s_locks_lower_in(17,18),
			in1                => s_in1(17,18),
			in2                => s_in2(17,18),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(18)
		);
	s_in1(17,18)            <= s_out1(18,18);
	s_in2(17,18)            <= s_out2(18,19);
	s_locks_lower_in(17,18) <= s_locks_lower_out(18,18);

		normal_cell_17_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,19),
			fetch              => s_fetch(17,19),
			data_in            => s_data_in(17,19),
			data_out           => s_data_out(17,19),
			out1               => s_out1(17,19),
			out2               => s_out2(17,19),
			lock_lower_row_out => s_locks_lower_out(17,19),
			lock_lower_row_in  => s_locks_lower_in(17,19),
			in1                => s_in1(17,19),
			in2                => s_in2(17,19),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(19)
		);
	s_in1(17,19)            <= s_out1(18,19);
	s_in2(17,19)            <= s_out2(18,20);
	s_locks_lower_in(17,19) <= s_locks_lower_out(18,19);

		normal_cell_17_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,20),
			fetch              => s_fetch(17,20),
			data_in            => s_data_in(17,20),
			data_out           => s_data_out(17,20),
			out1               => s_out1(17,20),
			out2               => s_out2(17,20),
			lock_lower_row_out => s_locks_lower_out(17,20),
			lock_lower_row_in  => s_locks_lower_in(17,20),
			in1                => s_in1(17,20),
			in2                => s_in2(17,20),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(20)
		);
	s_in1(17,20)            <= s_out1(18,20);
	s_in2(17,20)            <= s_out2(18,21);
	s_locks_lower_in(17,20) <= s_locks_lower_out(18,20);

		normal_cell_17_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,21),
			fetch              => s_fetch(17,21),
			data_in            => s_data_in(17,21),
			data_out           => s_data_out(17,21),
			out1               => s_out1(17,21),
			out2               => s_out2(17,21),
			lock_lower_row_out => s_locks_lower_out(17,21),
			lock_lower_row_in  => s_locks_lower_in(17,21),
			in1                => s_in1(17,21),
			in2                => s_in2(17,21),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(21)
		);
	s_in1(17,21)            <= s_out1(18,21);
	s_in2(17,21)            <= s_out2(18,22);
	s_locks_lower_in(17,21) <= s_locks_lower_out(18,21);

		normal_cell_17_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,22),
			fetch              => s_fetch(17,22),
			data_in            => s_data_in(17,22),
			data_out           => s_data_out(17,22),
			out1               => s_out1(17,22),
			out2               => s_out2(17,22),
			lock_lower_row_out => s_locks_lower_out(17,22),
			lock_lower_row_in  => s_locks_lower_in(17,22),
			in1                => s_in1(17,22),
			in2                => s_in2(17,22),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(22)
		);
	s_in1(17,22)            <= s_out1(18,22);
	s_in2(17,22)            <= s_out2(18,23);
	s_locks_lower_in(17,22) <= s_locks_lower_out(18,22);

		normal_cell_17_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,23),
			fetch              => s_fetch(17,23),
			data_in            => s_data_in(17,23),
			data_out           => s_data_out(17,23),
			out1               => s_out1(17,23),
			out2               => s_out2(17,23),
			lock_lower_row_out => s_locks_lower_out(17,23),
			lock_lower_row_in  => s_locks_lower_in(17,23),
			in1                => s_in1(17,23),
			in2                => s_in2(17,23),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(23)
		);
	s_in1(17,23)            <= s_out1(18,23);
	s_in2(17,23)            <= s_out2(18,24);
	s_locks_lower_in(17,23) <= s_locks_lower_out(18,23);

		normal_cell_17_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,24),
			fetch              => s_fetch(17,24),
			data_in            => s_data_in(17,24),
			data_out           => s_data_out(17,24),
			out1               => s_out1(17,24),
			out2               => s_out2(17,24),
			lock_lower_row_out => s_locks_lower_out(17,24),
			lock_lower_row_in  => s_locks_lower_in(17,24),
			in1                => s_in1(17,24),
			in2                => s_in2(17,24),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(24)
		);
	s_in1(17,24)            <= s_out1(18,24);
	s_in2(17,24)            <= s_out2(18,25);
	s_locks_lower_in(17,24) <= s_locks_lower_out(18,24);

		normal_cell_17_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,25),
			fetch              => s_fetch(17,25),
			data_in            => s_data_in(17,25),
			data_out           => s_data_out(17,25),
			out1               => s_out1(17,25),
			out2               => s_out2(17,25),
			lock_lower_row_out => s_locks_lower_out(17,25),
			lock_lower_row_in  => s_locks_lower_in(17,25),
			in1                => s_in1(17,25),
			in2                => s_in2(17,25),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(25)
		);
	s_in1(17,25)            <= s_out1(18,25);
	s_in2(17,25)            <= s_out2(18,26);
	s_locks_lower_in(17,25) <= s_locks_lower_out(18,25);

		normal_cell_17_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,26),
			fetch              => s_fetch(17,26),
			data_in            => s_data_in(17,26),
			data_out           => s_data_out(17,26),
			out1               => s_out1(17,26),
			out2               => s_out2(17,26),
			lock_lower_row_out => s_locks_lower_out(17,26),
			lock_lower_row_in  => s_locks_lower_in(17,26),
			in1                => s_in1(17,26),
			in2                => s_in2(17,26),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(26)
		);
	s_in1(17,26)            <= s_out1(18,26);
	s_in2(17,26)            <= s_out2(18,27);
	s_locks_lower_in(17,26) <= s_locks_lower_out(18,26);

		normal_cell_17_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,27),
			fetch              => s_fetch(17,27),
			data_in            => s_data_in(17,27),
			data_out           => s_data_out(17,27),
			out1               => s_out1(17,27),
			out2               => s_out2(17,27),
			lock_lower_row_out => s_locks_lower_out(17,27),
			lock_lower_row_in  => s_locks_lower_in(17,27),
			in1                => s_in1(17,27),
			in2                => s_in2(17,27),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(27)
		);
	s_in1(17,27)            <= s_out1(18,27);
	s_in2(17,27)            <= s_out2(18,28);
	s_locks_lower_in(17,27) <= s_locks_lower_out(18,27);

		normal_cell_17_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,28),
			fetch              => s_fetch(17,28),
			data_in            => s_data_in(17,28),
			data_out           => s_data_out(17,28),
			out1               => s_out1(17,28),
			out2               => s_out2(17,28),
			lock_lower_row_out => s_locks_lower_out(17,28),
			lock_lower_row_in  => s_locks_lower_in(17,28),
			in1                => s_in1(17,28),
			in2                => s_in2(17,28),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(28)
		);
	s_in1(17,28)            <= s_out1(18,28);
	s_in2(17,28)            <= s_out2(18,29);
	s_locks_lower_in(17,28) <= s_locks_lower_out(18,28);

		normal_cell_17_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,29),
			fetch              => s_fetch(17,29),
			data_in            => s_data_in(17,29),
			data_out           => s_data_out(17,29),
			out1               => s_out1(17,29),
			out2               => s_out2(17,29),
			lock_lower_row_out => s_locks_lower_out(17,29),
			lock_lower_row_in  => s_locks_lower_in(17,29),
			in1                => s_in1(17,29),
			in2                => s_in2(17,29),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(29)
		);
	s_in1(17,29)            <= s_out1(18,29);
	s_in2(17,29)            <= s_out2(18,30);
	s_locks_lower_in(17,29) <= s_locks_lower_out(18,29);

		normal_cell_17_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,30),
			fetch              => s_fetch(17,30),
			data_in            => s_data_in(17,30),
			data_out           => s_data_out(17,30),
			out1               => s_out1(17,30),
			out2               => s_out2(17,30),
			lock_lower_row_out => s_locks_lower_out(17,30),
			lock_lower_row_in  => s_locks_lower_in(17,30),
			in1                => s_in1(17,30),
			in2                => s_in2(17,30),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(30)
		);
	s_in1(17,30)            <= s_out1(18,30);
	s_in2(17,30)            <= s_out2(18,31);
	s_locks_lower_in(17,30) <= s_locks_lower_out(18,30);

		normal_cell_17_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,31),
			fetch              => s_fetch(17,31),
			data_in            => s_data_in(17,31),
			data_out           => s_data_out(17,31),
			out1               => s_out1(17,31),
			out2               => s_out2(17,31),
			lock_lower_row_out => s_locks_lower_out(17,31),
			lock_lower_row_in  => s_locks_lower_in(17,31),
			in1                => s_in1(17,31),
			in2                => s_in2(17,31),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(31)
		);
	s_in1(17,31)            <= s_out1(18,31);
	s_in2(17,31)            <= s_out2(18,32);
	s_locks_lower_in(17,31) <= s_locks_lower_out(18,31);

		normal_cell_17_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,32),
			fetch              => s_fetch(17,32),
			data_in            => s_data_in(17,32),
			data_out           => s_data_out(17,32),
			out1               => s_out1(17,32),
			out2               => s_out2(17,32),
			lock_lower_row_out => s_locks_lower_out(17,32),
			lock_lower_row_in  => s_locks_lower_in(17,32),
			in1                => s_in1(17,32),
			in2                => s_in2(17,32),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(32)
		);
	s_in1(17,32)            <= s_out1(18,32);
	s_in2(17,32)            <= s_out2(18,33);
	s_locks_lower_in(17,32) <= s_locks_lower_out(18,32);

		normal_cell_17_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,33),
			fetch              => s_fetch(17,33),
			data_in            => s_data_in(17,33),
			data_out           => s_data_out(17,33),
			out1               => s_out1(17,33),
			out2               => s_out2(17,33),
			lock_lower_row_out => s_locks_lower_out(17,33),
			lock_lower_row_in  => s_locks_lower_in(17,33),
			in1                => s_in1(17,33),
			in2                => s_in2(17,33),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(33)
		);
	s_in1(17,33)            <= s_out1(18,33);
	s_in2(17,33)            <= s_out2(18,34);
	s_locks_lower_in(17,33) <= s_locks_lower_out(18,33);

		normal_cell_17_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,34),
			fetch              => s_fetch(17,34),
			data_in            => s_data_in(17,34),
			data_out           => s_data_out(17,34),
			out1               => s_out1(17,34),
			out2               => s_out2(17,34),
			lock_lower_row_out => s_locks_lower_out(17,34),
			lock_lower_row_in  => s_locks_lower_in(17,34),
			in1                => s_in1(17,34),
			in2                => s_in2(17,34),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(34)
		);
	s_in1(17,34)            <= s_out1(18,34);
	s_in2(17,34)            <= s_out2(18,35);
	s_locks_lower_in(17,34) <= s_locks_lower_out(18,34);

		normal_cell_17_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,35),
			fetch              => s_fetch(17,35),
			data_in            => s_data_in(17,35),
			data_out           => s_data_out(17,35),
			out1               => s_out1(17,35),
			out2               => s_out2(17,35),
			lock_lower_row_out => s_locks_lower_out(17,35),
			lock_lower_row_in  => s_locks_lower_in(17,35),
			in1                => s_in1(17,35),
			in2                => s_in2(17,35),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(35)
		);
	s_in1(17,35)            <= s_out1(18,35);
	s_in2(17,35)            <= s_out2(18,36);
	s_locks_lower_in(17,35) <= s_locks_lower_out(18,35);

		normal_cell_17_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,36),
			fetch              => s_fetch(17,36),
			data_in            => s_data_in(17,36),
			data_out           => s_data_out(17,36),
			out1               => s_out1(17,36),
			out2               => s_out2(17,36),
			lock_lower_row_out => s_locks_lower_out(17,36),
			lock_lower_row_in  => s_locks_lower_in(17,36),
			in1                => s_in1(17,36),
			in2                => s_in2(17,36),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(36)
		);
	s_in1(17,36)            <= s_out1(18,36);
	s_in2(17,36)            <= s_out2(18,37);
	s_locks_lower_in(17,36) <= s_locks_lower_out(18,36);

		normal_cell_17_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,37),
			fetch              => s_fetch(17,37),
			data_in            => s_data_in(17,37),
			data_out           => s_data_out(17,37),
			out1               => s_out1(17,37),
			out2               => s_out2(17,37),
			lock_lower_row_out => s_locks_lower_out(17,37),
			lock_lower_row_in  => s_locks_lower_in(17,37),
			in1                => s_in1(17,37),
			in2                => s_in2(17,37),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(37)
		);
	s_in1(17,37)            <= s_out1(18,37);
	s_in2(17,37)            <= s_out2(18,38);
	s_locks_lower_in(17,37) <= s_locks_lower_out(18,37);

		normal_cell_17_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,38),
			fetch              => s_fetch(17,38),
			data_in            => s_data_in(17,38),
			data_out           => s_data_out(17,38),
			out1               => s_out1(17,38),
			out2               => s_out2(17,38),
			lock_lower_row_out => s_locks_lower_out(17,38),
			lock_lower_row_in  => s_locks_lower_in(17,38),
			in1                => s_in1(17,38),
			in2                => s_in2(17,38),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(38)
		);
	s_in1(17,38)            <= s_out1(18,38);
	s_in2(17,38)            <= s_out2(18,39);
	s_locks_lower_in(17,38) <= s_locks_lower_out(18,38);

		normal_cell_17_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,39),
			fetch              => s_fetch(17,39),
			data_in            => s_data_in(17,39),
			data_out           => s_data_out(17,39),
			out1               => s_out1(17,39),
			out2               => s_out2(17,39),
			lock_lower_row_out => s_locks_lower_out(17,39),
			lock_lower_row_in  => s_locks_lower_in(17,39),
			in1                => s_in1(17,39),
			in2                => s_in2(17,39),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(39)
		);
	s_in1(17,39)            <= s_out1(18,39);
	s_in2(17,39)            <= s_out2(18,40);
	s_locks_lower_in(17,39) <= s_locks_lower_out(18,39);

		normal_cell_17_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,40),
			fetch              => s_fetch(17,40),
			data_in            => s_data_in(17,40),
			data_out           => s_data_out(17,40),
			out1               => s_out1(17,40),
			out2               => s_out2(17,40),
			lock_lower_row_out => s_locks_lower_out(17,40),
			lock_lower_row_in  => s_locks_lower_in(17,40),
			in1                => s_in1(17,40),
			in2                => s_in2(17,40),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(40)
		);
	s_in1(17,40)            <= s_out1(18,40);
	s_in2(17,40)            <= s_out2(18,41);
	s_locks_lower_in(17,40) <= s_locks_lower_out(18,40);

		normal_cell_17_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,41),
			fetch              => s_fetch(17,41),
			data_in            => s_data_in(17,41),
			data_out           => s_data_out(17,41),
			out1               => s_out1(17,41),
			out2               => s_out2(17,41),
			lock_lower_row_out => s_locks_lower_out(17,41),
			lock_lower_row_in  => s_locks_lower_in(17,41),
			in1                => s_in1(17,41),
			in2                => s_in2(17,41),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(41)
		);
	s_in1(17,41)            <= s_out1(18,41);
	s_in2(17,41)            <= s_out2(18,42);
	s_locks_lower_in(17,41) <= s_locks_lower_out(18,41);

		normal_cell_17_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,42),
			fetch              => s_fetch(17,42),
			data_in            => s_data_in(17,42),
			data_out           => s_data_out(17,42),
			out1               => s_out1(17,42),
			out2               => s_out2(17,42),
			lock_lower_row_out => s_locks_lower_out(17,42),
			lock_lower_row_in  => s_locks_lower_in(17,42),
			in1                => s_in1(17,42),
			in2                => s_in2(17,42),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(42)
		);
	s_in1(17,42)            <= s_out1(18,42);
	s_in2(17,42)            <= s_out2(18,43);
	s_locks_lower_in(17,42) <= s_locks_lower_out(18,42);

		normal_cell_17_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,43),
			fetch              => s_fetch(17,43),
			data_in            => s_data_in(17,43),
			data_out           => s_data_out(17,43),
			out1               => s_out1(17,43),
			out2               => s_out2(17,43),
			lock_lower_row_out => s_locks_lower_out(17,43),
			lock_lower_row_in  => s_locks_lower_in(17,43),
			in1                => s_in1(17,43),
			in2                => s_in2(17,43),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(43)
		);
	s_in1(17,43)            <= s_out1(18,43);
	s_in2(17,43)            <= s_out2(18,44);
	s_locks_lower_in(17,43) <= s_locks_lower_out(18,43);

		normal_cell_17_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,44),
			fetch              => s_fetch(17,44),
			data_in            => s_data_in(17,44),
			data_out           => s_data_out(17,44),
			out1               => s_out1(17,44),
			out2               => s_out2(17,44),
			lock_lower_row_out => s_locks_lower_out(17,44),
			lock_lower_row_in  => s_locks_lower_in(17,44),
			in1                => s_in1(17,44),
			in2                => s_in2(17,44),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(44)
		);
	s_in1(17,44)            <= s_out1(18,44);
	s_in2(17,44)            <= s_out2(18,45);
	s_locks_lower_in(17,44) <= s_locks_lower_out(18,44);

		normal_cell_17_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,45),
			fetch              => s_fetch(17,45),
			data_in            => s_data_in(17,45),
			data_out           => s_data_out(17,45),
			out1               => s_out1(17,45),
			out2               => s_out2(17,45),
			lock_lower_row_out => s_locks_lower_out(17,45),
			lock_lower_row_in  => s_locks_lower_in(17,45),
			in1                => s_in1(17,45),
			in2                => s_in2(17,45),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(45)
		);
	s_in1(17,45)            <= s_out1(18,45);
	s_in2(17,45)            <= s_out2(18,46);
	s_locks_lower_in(17,45) <= s_locks_lower_out(18,45);

		normal_cell_17_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,46),
			fetch              => s_fetch(17,46),
			data_in            => s_data_in(17,46),
			data_out           => s_data_out(17,46),
			out1               => s_out1(17,46),
			out2               => s_out2(17,46),
			lock_lower_row_out => s_locks_lower_out(17,46),
			lock_lower_row_in  => s_locks_lower_in(17,46),
			in1                => s_in1(17,46),
			in2                => s_in2(17,46),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(46)
		);
	s_in1(17,46)            <= s_out1(18,46);
	s_in2(17,46)            <= s_out2(18,47);
	s_locks_lower_in(17,46) <= s_locks_lower_out(18,46);

		normal_cell_17_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,47),
			fetch              => s_fetch(17,47),
			data_in            => s_data_in(17,47),
			data_out           => s_data_out(17,47),
			out1               => s_out1(17,47),
			out2               => s_out2(17,47),
			lock_lower_row_out => s_locks_lower_out(17,47),
			lock_lower_row_in  => s_locks_lower_in(17,47),
			in1                => s_in1(17,47),
			in2                => s_in2(17,47),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(47)
		);
	s_in1(17,47)            <= s_out1(18,47);
	s_in2(17,47)            <= s_out2(18,48);
	s_locks_lower_in(17,47) <= s_locks_lower_out(18,47);

		normal_cell_17_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,48),
			fetch              => s_fetch(17,48),
			data_in            => s_data_in(17,48),
			data_out           => s_data_out(17,48),
			out1               => s_out1(17,48),
			out2               => s_out2(17,48),
			lock_lower_row_out => s_locks_lower_out(17,48),
			lock_lower_row_in  => s_locks_lower_in(17,48),
			in1                => s_in1(17,48),
			in2                => s_in2(17,48),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(48)
		);
	s_in1(17,48)            <= s_out1(18,48);
	s_in2(17,48)            <= s_out2(18,49);
	s_locks_lower_in(17,48) <= s_locks_lower_out(18,48);

		normal_cell_17_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,49),
			fetch              => s_fetch(17,49),
			data_in            => s_data_in(17,49),
			data_out           => s_data_out(17,49),
			out1               => s_out1(17,49),
			out2               => s_out2(17,49),
			lock_lower_row_out => s_locks_lower_out(17,49),
			lock_lower_row_in  => s_locks_lower_in(17,49),
			in1                => s_in1(17,49),
			in2                => s_in2(17,49),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(49)
		);
	s_in1(17,49)            <= s_out1(18,49);
	s_in2(17,49)            <= s_out2(18,50);
	s_locks_lower_in(17,49) <= s_locks_lower_out(18,49);

		normal_cell_17_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,50),
			fetch              => s_fetch(17,50),
			data_in            => s_data_in(17,50),
			data_out           => s_data_out(17,50),
			out1               => s_out1(17,50),
			out2               => s_out2(17,50),
			lock_lower_row_out => s_locks_lower_out(17,50),
			lock_lower_row_in  => s_locks_lower_in(17,50),
			in1                => s_in1(17,50),
			in2                => s_in2(17,50),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(50)
		);
	s_in1(17,50)            <= s_out1(18,50);
	s_in2(17,50)            <= s_out2(18,51);
	s_locks_lower_in(17,50) <= s_locks_lower_out(18,50);

		normal_cell_17_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,51),
			fetch              => s_fetch(17,51),
			data_in            => s_data_in(17,51),
			data_out           => s_data_out(17,51),
			out1               => s_out1(17,51),
			out2               => s_out2(17,51),
			lock_lower_row_out => s_locks_lower_out(17,51),
			lock_lower_row_in  => s_locks_lower_in(17,51),
			in1                => s_in1(17,51),
			in2                => s_in2(17,51),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(51)
		);
	s_in1(17,51)            <= s_out1(18,51);
	s_in2(17,51)            <= s_out2(18,52);
	s_locks_lower_in(17,51) <= s_locks_lower_out(18,51);

		normal_cell_17_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,52),
			fetch              => s_fetch(17,52),
			data_in            => s_data_in(17,52),
			data_out           => s_data_out(17,52),
			out1               => s_out1(17,52),
			out2               => s_out2(17,52),
			lock_lower_row_out => s_locks_lower_out(17,52),
			lock_lower_row_in  => s_locks_lower_in(17,52),
			in1                => s_in1(17,52),
			in2                => s_in2(17,52),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(52)
		);
	s_in1(17,52)            <= s_out1(18,52);
	s_in2(17,52)            <= s_out2(18,53);
	s_locks_lower_in(17,52) <= s_locks_lower_out(18,52);

		normal_cell_17_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,53),
			fetch              => s_fetch(17,53),
			data_in            => s_data_in(17,53),
			data_out           => s_data_out(17,53),
			out1               => s_out1(17,53),
			out2               => s_out2(17,53),
			lock_lower_row_out => s_locks_lower_out(17,53),
			lock_lower_row_in  => s_locks_lower_in(17,53),
			in1                => s_in1(17,53),
			in2                => s_in2(17,53),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(53)
		);
	s_in1(17,53)            <= s_out1(18,53);
	s_in2(17,53)            <= s_out2(18,54);
	s_locks_lower_in(17,53) <= s_locks_lower_out(18,53);

		normal_cell_17_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,54),
			fetch              => s_fetch(17,54),
			data_in            => s_data_in(17,54),
			data_out           => s_data_out(17,54),
			out1               => s_out1(17,54),
			out2               => s_out2(17,54),
			lock_lower_row_out => s_locks_lower_out(17,54),
			lock_lower_row_in  => s_locks_lower_in(17,54),
			in1                => s_in1(17,54),
			in2                => s_in2(17,54),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(54)
		);
	s_in1(17,54)            <= s_out1(18,54);
	s_in2(17,54)            <= s_out2(18,55);
	s_locks_lower_in(17,54) <= s_locks_lower_out(18,54);

		normal_cell_17_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,55),
			fetch              => s_fetch(17,55),
			data_in            => s_data_in(17,55),
			data_out           => s_data_out(17,55),
			out1               => s_out1(17,55),
			out2               => s_out2(17,55),
			lock_lower_row_out => s_locks_lower_out(17,55),
			lock_lower_row_in  => s_locks_lower_in(17,55),
			in1                => s_in1(17,55),
			in2                => s_in2(17,55),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(55)
		);
	s_in1(17,55)            <= s_out1(18,55);
	s_in2(17,55)            <= s_out2(18,56);
	s_locks_lower_in(17,55) <= s_locks_lower_out(18,55);

		normal_cell_17_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,56),
			fetch              => s_fetch(17,56),
			data_in            => s_data_in(17,56),
			data_out           => s_data_out(17,56),
			out1               => s_out1(17,56),
			out2               => s_out2(17,56),
			lock_lower_row_out => s_locks_lower_out(17,56),
			lock_lower_row_in  => s_locks_lower_in(17,56),
			in1                => s_in1(17,56),
			in2                => s_in2(17,56),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(56)
		);
	s_in1(17,56)            <= s_out1(18,56);
	s_in2(17,56)            <= s_out2(18,57);
	s_locks_lower_in(17,56) <= s_locks_lower_out(18,56);

		normal_cell_17_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,57),
			fetch              => s_fetch(17,57),
			data_in            => s_data_in(17,57),
			data_out           => s_data_out(17,57),
			out1               => s_out1(17,57),
			out2               => s_out2(17,57),
			lock_lower_row_out => s_locks_lower_out(17,57),
			lock_lower_row_in  => s_locks_lower_in(17,57),
			in1                => s_in1(17,57),
			in2                => s_in2(17,57),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(57)
		);
	s_in1(17,57)            <= s_out1(18,57);
	s_in2(17,57)            <= s_out2(18,58);
	s_locks_lower_in(17,57) <= s_locks_lower_out(18,57);

		normal_cell_17_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,58),
			fetch              => s_fetch(17,58),
			data_in            => s_data_in(17,58),
			data_out           => s_data_out(17,58),
			out1               => s_out1(17,58),
			out2               => s_out2(17,58),
			lock_lower_row_out => s_locks_lower_out(17,58),
			lock_lower_row_in  => s_locks_lower_in(17,58),
			in1                => s_in1(17,58),
			in2                => s_in2(17,58),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(58)
		);
	s_in1(17,58)            <= s_out1(18,58);
	s_in2(17,58)            <= s_out2(18,59);
	s_locks_lower_in(17,58) <= s_locks_lower_out(18,58);

		normal_cell_17_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,59),
			fetch              => s_fetch(17,59),
			data_in            => s_data_in(17,59),
			data_out           => s_data_out(17,59),
			out1               => s_out1(17,59),
			out2               => s_out2(17,59),
			lock_lower_row_out => s_locks_lower_out(17,59),
			lock_lower_row_in  => s_locks_lower_in(17,59),
			in1                => s_in1(17,59),
			in2                => s_in2(17,59),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(59)
		);
	s_in1(17,59)            <= s_out1(18,59);
	s_in2(17,59)            <= s_out2(18,60);
	s_locks_lower_in(17,59) <= s_locks_lower_out(18,59);

		last_col_cell_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(17,60),
			fetch              => s_fetch(17,60),
			data_in            => s_data_in(17,60),
			data_out           => s_data_out(17,60),
			out1               => s_out1(17,60),
			out2               => s_out2(17,60),
			lock_lower_row_out => s_locks_lower_out(17,60),
			lock_lower_row_in  => s_locks_lower_in(17,60),
			in1                => s_in1(17,60),
			in2                => (others => '0'),
			lock_row           => s_locks(17),
			piv_found          => s_piv_found,
			row_data           => s_row_data(17),
			col_data           => s_col_data(60)
		);
	s_in1(17,60)            <= s_out1(18,60);
	s_locks_lower_in(17,60) <= s_locks_lower_out(18,60);

		normal_cell_18_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,1),
			fetch              => s_fetch(18,1),
			data_in            => s_data_in(18,1),
			data_out           => s_data_out(18,1),
			out1               => s_out1(18,1),
			out2               => s_out2(18,1),
			lock_lower_row_out => s_locks_lower_out(18,1),
			lock_lower_row_in  => s_locks_lower_in(18,1),
			in1                => s_in1(18,1),
			in2                => s_in2(18,1),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(1)
		);
	s_in1(18,1)            <= s_out1(19,1);
	s_in2(18,1)            <= s_out2(19,2);
	s_locks_lower_in(18,1) <= s_locks_lower_out(19,1);

		normal_cell_18_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,2),
			fetch              => s_fetch(18,2),
			data_in            => s_data_in(18,2),
			data_out           => s_data_out(18,2),
			out1               => s_out1(18,2),
			out2               => s_out2(18,2),
			lock_lower_row_out => s_locks_lower_out(18,2),
			lock_lower_row_in  => s_locks_lower_in(18,2),
			in1                => s_in1(18,2),
			in2                => s_in2(18,2),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(2)
		);
	s_in1(18,2)            <= s_out1(19,2);
	s_in2(18,2)            <= s_out2(19,3);
	s_locks_lower_in(18,2) <= s_locks_lower_out(19,2);

		normal_cell_18_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,3),
			fetch              => s_fetch(18,3),
			data_in            => s_data_in(18,3),
			data_out           => s_data_out(18,3),
			out1               => s_out1(18,3),
			out2               => s_out2(18,3),
			lock_lower_row_out => s_locks_lower_out(18,3),
			lock_lower_row_in  => s_locks_lower_in(18,3),
			in1                => s_in1(18,3),
			in2                => s_in2(18,3),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(3)
		);
	s_in1(18,3)            <= s_out1(19,3);
	s_in2(18,3)            <= s_out2(19,4);
	s_locks_lower_in(18,3) <= s_locks_lower_out(19,3);

		normal_cell_18_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,4),
			fetch              => s_fetch(18,4),
			data_in            => s_data_in(18,4),
			data_out           => s_data_out(18,4),
			out1               => s_out1(18,4),
			out2               => s_out2(18,4),
			lock_lower_row_out => s_locks_lower_out(18,4),
			lock_lower_row_in  => s_locks_lower_in(18,4),
			in1                => s_in1(18,4),
			in2                => s_in2(18,4),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(4)
		);
	s_in1(18,4)            <= s_out1(19,4);
	s_in2(18,4)            <= s_out2(19,5);
	s_locks_lower_in(18,4) <= s_locks_lower_out(19,4);

		normal_cell_18_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,5),
			fetch              => s_fetch(18,5),
			data_in            => s_data_in(18,5),
			data_out           => s_data_out(18,5),
			out1               => s_out1(18,5),
			out2               => s_out2(18,5),
			lock_lower_row_out => s_locks_lower_out(18,5),
			lock_lower_row_in  => s_locks_lower_in(18,5),
			in1                => s_in1(18,5),
			in2                => s_in2(18,5),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(5)
		);
	s_in1(18,5)            <= s_out1(19,5);
	s_in2(18,5)            <= s_out2(19,6);
	s_locks_lower_in(18,5) <= s_locks_lower_out(19,5);

		normal_cell_18_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,6),
			fetch              => s_fetch(18,6),
			data_in            => s_data_in(18,6),
			data_out           => s_data_out(18,6),
			out1               => s_out1(18,6),
			out2               => s_out2(18,6),
			lock_lower_row_out => s_locks_lower_out(18,6),
			lock_lower_row_in  => s_locks_lower_in(18,6),
			in1                => s_in1(18,6),
			in2                => s_in2(18,6),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(6)
		);
	s_in1(18,6)            <= s_out1(19,6);
	s_in2(18,6)            <= s_out2(19,7);
	s_locks_lower_in(18,6) <= s_locks_lower_out(19,6);

		normal_cell_18_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,7),
			fetch              => s_fetch(18,7),
			data_in            => s_data_in(18,7),
			data_out           => s_data_out(18,7),
			out1               => s_out1(18,7),
			out2               => s_out2(18,7),
			lock_lower_row_out => s_locks_lower_out(18,7),
			lock_lower_row_in  => s_locks_lower_in(18,7),
			in1                => s_in1(18,7),
			in2                => s_in2(18,7),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(7)
		);
	s_in1(18,7)            <= s_out1(19,7);
	s_in2(18,7)            <= s_out2(19,8);
	s_locks_lower_in(18,7) <= s_locks_lower_out(19,7);

		normal_cell_18_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,8),
			fetch              => s_fetch(18,8),
			data_in            => s_data_in(18,8),
			data_out           => s_data_out(18,8),
			out1               => s_out1(18,8),
			out2               => s_out2(18,8),
			lock_lower_row_out => s_locks_lower_out(18,8),
			lock_lower_row_in  => s_locks_lower_in(18,8),
			in1                => s_in1(18,8),
			in2                => s_in2(18,8),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(8)
		);
	s_in1(18,8)            <= s_out1(19,8);
	s_in2(18,8)            <= s_out2(19,9);
	s_locks_lower_in(18,8) <= s_locks_lower_out(19,8);

		normal_cell_18_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,9),
			fetch              => s_fetch(18,9),
			data_in            => s_data_in(18,9),
			data_out           => s_data_out(18,9),
			out1               => s_out1(18,9),
			out2               => s_out2(18,9),
			lock_lower_row_out => s_locks_lower_out(18,9),
			lock_lower_row_in  => s_locks_lower_in(18,9),
			in1                => s_in1(18,9),
			in2                => s_in2(18,9),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(9)
		);
	s_in1(18,9)            <= s_out1(19,9);
	s_in2(18,9)            <= s_out2(19,10);
	s_locks_lower_in(18,9) <= s_locks_lower_out(19,9);

		normal_cell_18_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,10),
			fetch              => s_fetch(18,10),
			data_in            => s_data_in(18,10),
			data_out           => s_data_out(18,10),
			out1               => s_out1(18,10),
			out2               => s_out2(18,10),
			lock_lower_row_out => s_locks_lower_out(18,10),
			lock_lower_row_in  => s_locks_lower_in(18,10),
			in1                => s_in1(18,10),
			in2                => s_in2(18,10),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(10)
		);
	s_in1(18,10)            <= s_out1(19,10);
	s_in2(18,10)            <= s_out2(19,11);
	s_locks_lower_in(18,10) <= s_locks_lower_out(19,10);

		normal_cell_18_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,11),
			fetch              => s_fetch(18,11),
			data_in            => s_data_in(18,11),
			data_out           => s_data_out(18,11),
			out1               => s_out1(18,11),
			out2               => s_out2(18,11),
			lock_lower_row_out => s_locks_lower_out(18,11),
			lock_lower_row_in  => s_locks_lower_in(18,11),
			in1                => s_in1(18,11),
			in2                => s_in2(18,11),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(11)
		);
	s_in1(18,11)            <= s_out1(19,11);
	s_in2(18,11)            <= s_out2(19,12);
	s_locks_lower_in(18,11) <= s_locks_lower_out(19,11);

		normal_cell_18_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,12),
			fetch              => s_fetch(18,12),
			data_in            => s_data_in(18,12),
			data_out           => s_data_out(18,12),
			out1               => s_out1(18,12),
			out2               => s_out2(18,12),
			lock_lower_row_out => s_locks_lower_out(18,12),
			lock_lower_row_in  => s_locks_lower_in(18,12),
			in1                => s_in1(18,12),
			in2                => s_in2(18,12),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(12)
		);
	s_in1(18,12)            <= s_out1(19,12);
	s_in2(18,12)            <= s_out2(19,13);
	s_locks_lower_in(18,12) <= s_locks_lower_out(19,12);

		normal_cell_18_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,13),
			fetch              => s_fetch(18,13),
			data_in            => s_data_in(18,13),
			data_out           => s_data_out(18,13),
			out1               => s_out1(18,13),
			out2               => s_out2(18,13),
			lock_lower_row_out => s_locks_lower_out(18,13),
			lock_lower_row_in  => s_locks_lower_in(18,13),
			in1                => s_in1(18,13),
			in2                => s_in2(18,13),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(13)
		);
	s_in1(18,13)            <= s_out1(19,13);
	s_in2(18,13)            <= s_out2(19,14);
	s_locks_lower_in(18,13) <= s_locks_lower_out(19,13);

		normal_cell_18_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,14),
			fetch              => s_fetch(18,14),
			data_in            => s_data_in(18,14),
			data_out           => s_data_out(18,14),
			out1               => s_out1(18,14),
			out2               => s_out2(18,14),
			lock_lower_row_out => s_locks_lower_out(18,14),
			lock_lower_row_in  => s_locks_lower_in(18,14),
			in1                => s_in1(18,14),
			in2                => s_in2(18,14),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(14)
		);
	s_in1(18,14)            <= s_out1(19,14);
	s_in2(18,14)            <= s_out2(19,15);
	s_locks_lower_in(18,14) <= s_locks_lower_out(19,14);

		normal_cell_18_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,15),
			fetch              => s_fetch(18,15),
			data_in            => s_data_in(18,15),
			data_out           => s_data_out(18,15),
			out1               => s_out1(18,15),
			out2               => s_out2(18,15),
			lock_lower_row_out => s_locks_lower_out(18,15),
			lock_lower_row_in  => s_locks_lower_in(18,15),
			in1                => s_in1(18,15),
			in2                => s_in2(18,15),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(15)
		);
	s_in1(18,15)            <= s_out1(19,15);
	s_in2(18,15)            <= s_out2(19,16);
	s_locks_lower_in(18,15) <= s_locks_lower_out(19,15);

		normal_cell_18_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,16),
			fetch              => s_fetch(18,16),
			data_in            => s_data_in(18,16),
			data_out           => s_data_out(18,16),
			out1               => s_out1(18,16),
			out2               => s_out2(18,16),
			lock_lower_row_out => s_locks_lower_out(18,16),
			lock_lower_row_in  => s_locks_lower_in(18,16),
			in1                => s_in1(18,16),
			in2                => s_in2(18,16),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(16)
		);
	s_in1(18,16)            <= s_out1(19,16);
	s_in2(18,16)            <= s_out2(19,17);
	s_locks_lower_in(18,16) <= s_locks_lower_out(19,16);

		normal_cell_18_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,17),
			fetch              => s_fetch(18,17),
			data_in            => s_data_in(18,17),
			data_out           => s_data_out(18,17),
			out1               => s_out1(18,17),
			out2               => s_out2(18,17),
			lock_lower_row_out => s_locks_lower_out(18,17),
			lock_lower_row_in  => s_locks_lower_in(18,17),
			in1                => s_in1(18,17),
			in2                => s_in2(18,17),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(17)
		);
	s_in1(18,17)            <= s_out1(19,17);
	s_in2(18,17)            <= s_out2(19,18);
	s_locks_lower_in(18,17) <= s_locks_lower_out(19,17);

		normal_cell_18_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,18),
			fetch              => s_fetch(18,18),
			data_in            => s_data_in(18,18),
			data_out           => s_data_out(18,18),
			out1               => s_out1(18,18),
			out2               => s_out2(18,18),
			lock_lower_row_out => s_locks_lower_out(18,18),
			lock_lower_row_in  => s_locks_lower_in(18,18),
			in1                => s_in1(18,18),
			in2                => s_in2(18,18),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(18)
		);
	s_in1(18,18)            <= s_out1(19,18);
	s_in2(18,18)            <= s_out2(19,19);
	s_locks_lower_in(18,18) <= s_locks_lower_out(19,18);

		normal_cell_18_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,19),
			fetch              => s_fetch(18,19),
			data_in            => s_data_in(18,19),
			data_out           => s_data_out(18,19),
			out1               => s_out1(18,19),
			out2               => s_out2(18,19),
			lock_lower_row_out => s_locks_lower_out(18,19),
			lock_lower_row_in  => s_locks_lower_in(18,19),
			in1                => s_in1(18,19),
			in2                => s_in2(18,19),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(19)
		);
	s_in1(18,19)            <= s_out1(19,19);
	s_in2(18,19)            <= s_out2(19,20);
	s_locks_lower_in(18,19) <= s_locks_lower_out(19,19);

		normal_cell_18_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,20),
			fetch              => s_fetch(18,20),
			data_in            => s_data_in(18,20),
			data_out           => s_data_out(18,20),
			out1               => s_out1(18,20),
			out2               => s_out2(18,20),
			lock_lower_row_out => s_locks_lower_out(18,20),
			lock_lower_row_in  => s_locks_lower_in(18,20),
			in1                => s_in1(18,20),
			in2                => s_in2(18,20),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(20)
		);
	s_in1(18,20)            <= s_out1(19,20);
	s_in2(18,20)            <= s_out2(19,21);
	s_locks_lower_in(18,20) <= s_locks_lower_out(19,20);

		normal_cell_18_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,21),
			fetch              => s_fetch(18,21),
			data_in            => s_data_in(18,21),
			data_out           => s_data_out(18,21),
			out1               => s_out1(18,21),
			out2               => s_out2(18,21),
			lock_lower_row_out => s_locks_lower_out(18,21),
			lock_lower_row_in  => s_locks_lower_in(18,21),
			in1                => s_in1(18,21),
			in2                => s_in2(18,21),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(21)
		);
	s_in1(18,21)            <= s_out1(19,21);
	s_in2(18,21)            <= s_out2(19,22);
	s_locks_lower_in(18,21) <= s_locks_lower_out(19,21);

		normal_cell_18_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,22),
			fetch              => s_fetch(18,22),
			data_in            => s_data_in(18,22),
			data_out           => s_data_out(18,22),
			out1               => s_out1(18,22),
			out2               => s_out2(18,22),
			lock_lower_row_out => s_locks_lower_out(18,22),
			lock_lower_row_in  => s_locks_lower_in(18,22),
			in1                => s_in1(18,22),
			in2                => s_in2(18,22),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(22)
		);
	s_in1(18,22)            <= s_out1(19,22);
	s_in2(18,22)            <= s_out2(19,23);
	s_locks_lower_in(18,22) <= s_locks_lower_out(19,22);

		normal_cell_18_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,23),
			fetch              => s_fetch(18,23),
			data_in            => s_data_in(18,23),
			data_out           => s_data_out(18,23),
			out1               => s_out1(18,23),
			out2               => s_out2(18,23),
			lock_lower_row_out => s_locks_lower_out(18,23),
			lock_lower_row_in  => s_locks_lower_in(18,23),
			in1                => s_in1(18,23),
			in2                => s_in2(18,23),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(23)
		);
	s_in1(18,23)            <= s_out1(19,23);
	s_in2(18,23)            <= s_out2(19,24);
	s_locks_lower_in(18,23) <= s_locks_lower_out(19,23);

		normal_cell_18_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,24),
			fetch              => s_fetch(18,24),
			data_in            => s_data_in(18,24),
			data_out           => s_data_out(18,24),
			out1               => s_out1(18,24),
			out2               => s_out2(18,24),
			lock_lower_row_out => s_locks_lower_out(18,24),
			lock_lower_row_in  => s_locks_lower_in(18,24),
			in1                => s_in1(18,24),
			in2                => s_in2(18,24),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(24)
		);
	s_in1(18,24)            <= s_out1(19,24);
	s_in2(18,24)            <= s_out2(19,25);
	s_locks_lower_in(18,24) <= s_locks_lower_out(19,24);

		normal_cell_18_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,25),
			fetch              => s_fetch(18,25),
			data_in            => s_data_in(18,25),
			data_out           => s_data_out(18,25),
			out1               => s_out1(18,25),
			out2               => s_out2(18,25),
			lock_lower_row_out => s_locks_lower_out(18,25),
			lock_lower_row_in  => s_locks_lower_in(18,25),
			in1                => s_in1(18,25),
			in2                => s_in2(18,25),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(25)
		);
	s_in1(18,25)            <= s_out1(19,25);
	s_in2(18,25)            <= s_out2(19,26);
	s_locks_lower_in(18,25) <= s_locks_lower_out(19,25);

		normal_cell_18_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,26),
			fetch              => s_fetch(18,26),
			data_in            => s_data_in(18,26),
			data_out           => s_data_out(18,26),
			out1               => s_out1(18,26),
			out2               => s_out2(18,26),
			lock_lower_row_out => s_locks_lower_out(18,26),
			lock_lower_row_in  => s_locks_lower_in(18,26),
			in1                => s_in1(18,26),
			in2                => s_in2(18,26),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(26)
		);
	s_in1(18,26)            <= s_out1(19,26);
	s_in2(18,26)            <= s_out2(19,27);
	s_locks_lower_in(18,26) <= s_locks_lower_out(19,26);

		normal_cell_18_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,27),
			fetch              => s_fetch(18,27),
			data_in            => s_data_in(18,27),
			data_out           => s_data_out(18,27),
			out1               => s_out1(18,27),
			out2               => s_out2(18,27),
			lock_lower_row_out => s_locks_lower_out(18,27),
			lock_lower_row_in  => s_locks_lower_in(18,27),
			in1                => s_in1(18,27),
			in2                => s_in2(18,27),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(27)
		);
	s_in1(18,27)            <= s_out1(19,27);
	s_in2(18,27)            <= s_out2(19,28);
	s_locks_lower_in(18,27) <= s_locks_lower_out(19,27);

		normal_cell_18_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,28),
			fetch              => s_fetch(18,28),
			data_in            => s_data_in(18,28),
			data_out           => s_data_out(18,28),
			out1               => s_out1(18,28),
			out2               => s_out2(18,28),
			lock_lower_row_out => s_locks_lower_out(18,28),
			lock_lower_row_in  => s_locks_lower_in(18,28),
			in1                => s_in1(18,28),
			in2                => s_in2(18,28),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(28)
		);
	s_in1(18,28)            <= s_out1(19,28);
	s_in2(18,28)            <= s_out2(19,29);
	s_locks_lower_in(18,28) <= s_locks_lower_out(19,28);

		normal_cell_18_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,29),
			fetch              => s_fetch(18,29),
			data_in            => s_data_in(18,29),
			data_out           => s_data_out(18,29),
			out1               => s_out1(18,29),
			out2               => s_out2(18,29),
			lock_lower_row_out => s_locks_lower_out(18,29),
			lock_lower_row_in  => s_locks_lower_in(18,29),
			in1                => s_in1(18,29),
			in2                => s_in2(18,29),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(29)
		);
	s_in1(18,29)            <= s_out1(19,29);
	s_in2(18,29)            <= s_out2(19,30);
	s_locks_lower_in(18,29) <= s_locks_lower_out(19,29);

		normal_cell_18_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,30),
			fetch              => s_fetch(18,30),
			data_in            => s_data_in(18,30),
			data_out           => s_data_out(18,30),
			out1               => s_out1(18,30),
			out2               => s_out2(18,30),
			lock_lower_row_out => s_locks_lower_out(18,30),
			lock_lower_row_in  => s_locks_lower_in(18,30),
			in1                => s_in1(18,30),
			in2                => s_in2(18,30),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(30)
		);
	s_in1(18,30)            <= s_out1(19,30);
	s_in2(18,30)            <= s_out2(19,31);
	s_locks_lower_in(18,30) <= s_locks_lower_out(19,30);

		normal_cell_18_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,31),
			fetch              => s_fetch(18,31),
			data_in            => s_data_in(18,31),
			data_out           => s_data_out(18,31),
			out1               => s_out1(18,31),
			out2               => s_out2(18,31),
			lock_lower_row_out => s_locks_lower_out(18,31),
			lock_lower_row_in  => s_locks_lower_in(18,31),
			in1                => s_in1(18,31),
			in2                => s_in2(18,31),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(31)
		);
	s_in1(18,31)            <= s_out1(19,31);
	s_in2(18,31)            <= s_out2(19,32);
	s_locks_lower_in(18,31) <= s_locks_lower_out(19,31);

		normal_cell_18_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,32),
			fetch              => s_fetch(18,32),
			data_in            => s_data_in(18,32),
			data_out           => s_data_out(18,32),
			out1               => s_out1(18,32),
			out2               => s_out2(18,32),
			lock_lower_row_out => s_locks_lower_out(18,32),
			lock_lower_row_in  => s_locks_lower_in(18,32),
			in1                => s_in1(18,32),
			in2                => s_in2(18,32),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(32)
		);
	s_in1(18,32)            <= s_out1(19,32);
	s_in2(18,32)            <= s_out2(19,33);
	s_locks_lower_in(18,32) <= s_locks_lower_out(19,32);

		normal_cell_18_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,33),
			fetch              => s_fetch(18,33),
			data_in            => s_data_in(18,33),
			data_out           => s_data_out(18,33),
			out1               => s_out1(18,33),
			out2               => s_out2(18,33),
			lock_lower_row_out => s_locks_lower_out(18,33),
			lock_lower_row_in  => s_locks_lower_in(18,33),
			in1                => s_in1(18,33),
			in2                => s_in2(18,33),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(33)
		);
	s_in1(18,33)            <= s_out1(19,33);
	s_in2(18,33)            <= s_out2(19,34);
	s_locks_lower_in(18,33) <= s_locks_lower_out(19,33);

		normal_cell_18_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,34),
			fetch              => s_fetch(18,34),
			data_in            => s_data_in(18,34),
			data_out           => s_data_out(18,34),
			out1               => s_out1(18,34),
			out2               => s_out2(18,34),
			lock_lower_row_out => s_locks_lower_out(18,34),
			lock_lower_row_in  => s_locks_lower_in(18,34),
			in1                => s_in1(18,34),
			in2                => s_in2(18,34),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(34)
		);
	s_in1(18,34)            <= s_out1(19,34);
	s_in2(18,34)            <= s_out2(19,35);
	s_locks_lower_in(18,34) <= s_locks_lower_out(19,34);

		normal_cell_18_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,35),
			fetch              => s_fetch(18,35),
			data_in            => s_data_in(18,35),
			data_out           => s_data_out(18,35),
			out1               => s_out1(18,35),
			out2               => s_out2(18,35),
			lock_lower_row_out => s_locks_lower_out(18,35),
			lock_lower_row_in  => s_locks_lower_in(18,35),
			in1                => s_in1(18,35),
			in2                => s_in2(18,35),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(35)
		);
	s_in1(18,35)            <= s_out1(19,35);
	s_in2(18,35)            <= s_out2(19,36);
	s_locks_lower_in(18,35) <= s_locks_lower_out(19,35);

		normal_cell_18_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,36),
			fetch              => s_fetch(18,36),
			data_in            => s_data_in(18,36),
			data_out           => s_data_out(18,36),
			out1               => s_out1(18,36),
			out2               => s_out2(18,36),
			lock_lower_row_out => s_locks_lower_out(18,36),
			lock_lower_row_in  => s_locks_lower_in(18,36),
			in1                => s_in1(18,36),
			in2                => s_in2(18,36),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(36)
		);
	s_in1(18,36)            <= s_out1(19,36);
	s_in2(18,36)            <= s_out2(19,37);
	s_locks_lower_in(18,36) <= s_locks_lower_out(19,36);

		normal_cell_18_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,37),
			fetch              => s_fetch(18,37),
			data_in            => s_data_in(18,37),
			data_out           => s_data_out(18,37),
			out1               => s_out1(18,37),
			out2               => s_out2(18,37),
			lock_lower_row_out => s_locks_lower_out(18,37),
			lock_lower_row_in  => s_locks_lower_in(18,37),
			in1                => s_in1(18,37),
			in2                => s_in2(18,37),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(37)
		);
	s_in1(18,37)            <= s_out1(19,37);
	s_in2(18,37)            <= s_out2(19,38);
	s_locks_lower_in(18,37) <= s_locks_lower_out(19,37);

		normal_cell_18_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,38),
			fetch              => s_fetch(18,38),
			data_in            => s_data_in(18,38),
			data_out           => s_data_out(18,38),
			out1               => s_out1(18,38),
			out2               => s_out2(18,38),
			lock_lower_row_out => s_locks_lower_out(18,38),
			lock_lower_row_in  => s_locks_lower_in(18,38),
			in1                => s_in1(18,38),
			in2                => s_in2(18,38),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(38)
		);
	s_in1(18,38)            <= s_out1(19,38);
	s_in2(18,38)            <= s_out2(19,39);
	s_locks_lower_in(18,38) <= s_locks_lower_out(19,38);

		normal_cell_18_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,39),
			fetch              => s_fetch(18,39),
			data_in            => s_data_in(18,39),
			data_out           => s_data_out(18,39),
			out1               => s_out1(18,39),
			out2               => s_out2(18,39),
			lock_lower_row_out => s_locks_lower_out(18,39),
			lock_lower_row_in  => s_locks_lower_in(18,39),
			in1                => s_in1(18,39),
			in2                => s_in2(18,39),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(39)
		);
	s_in1(18,39)            <= s_out1(19,39);
	s_in2(18,39)            <= s_out2(19,40);
	s_locks_lower_in(18,39) <= s_locks_lower_out(19,39);

		normal_cell_18_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,40),
			fetch              => s_fetch(18,40),
			data_in            => s_data_in(18,40),
			data_out           => s_data_out(18,40),
			out1               => s_out1(18,40),
			out2               => s_out2(18,40),
			lock_lower_row_out => s_locks_lower_out(18,40),
			lock_lower_row_in  => s_locks_lower_in(18,40),
			in1                => s_in1(18,40),
			in2                => s_in2(18,40),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(40)
		);
	s_in1(18,40)            <= s_out1(19,40);
	s_in2(18,40)            <= s_out2(19,41);
	s_locks_lower_in(18,40) <= s_locks_lower_out(19,40);

		normal_cell_18_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,41),
			fetch              => s_fetch(18,41),
			data_in            => s_data_in(18,41),
			data_out           => s_data_out(18,41),
			out1               => s_out1(18,41),
			out2               => s_out2(18,41),
			lock_lower_row_out => s_locks_lower_out(18,41),
			lock_lower_row_in  => s_locks_lower_in(18,41),
			in1                => s_in1(18,41),
			in2                => s_in2(18,41),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(41)
		);
	s_in1(18,41)            <= s_out1(19,41);
	s_in2(18,41)            <= s_out2(19,42);
	s_locks_lower_in(18,41) <= s_locks_lower_out(19,41);

		normal_cell_18_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,42),
			fetch              => s_fetch(18,42),
			data_in            => s_data_in(18,42),
			data_out           => s_data_out(18,42),
			out1               => s_out1(18,42),
			out2               => s_out2(18,42),
			lock_lower_row_out => s_locks_lower_out(18,42),
			lock_lower_row_in  => s_locks_lower_in(18,42),
			in1                => s_in1(18,42),
			in2                => s_in2(18,42),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(42)
		);
	s_in1(18,42)            <= s_out1(19,42);
	s_in2(18,42)            <= s_out2(19,43);
	s_locks_lower_in(18,42) <= s_locks_lower_out(19,42);

		normal_cell_18_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,43),
			fetch              => s_fetch(18,43),
			data_in            => s_data_in(18,43),
			data_out           => s_data_out(18,43),
			out1               => s_out1(18,43),
			out2               => s_out2(18,43),
			lock_lower_row_out => s_locks_lower_out(18,43),
			lock_lower_row_in  => s_locks_lower_in(18,43),
			in1                => s_in1(18,43),
			in2                => s_in2(18,43),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(43)
		);
	s_in1(18,43)            <= s_out1(19,43);
	s_in2(18,43)            <= s_out2(19,44);
	s_locks_lower_in(18,43) <= s_locks_lower_out(19,43);

		normal_cell_18_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,44),
			fetch              => s_fetch(18,44),
			data_in            => s_data_in(18,44),
			data_out           => s_data_out(18,44),
			out1               => s_out1(18,44),
			out2               => s_out2(18,44),
			lock_lower_row_out => s_locks_lower_out(18,44),
			lock_lower_row_in  => s_locks_lower_in(18,44),
			in1                => s_in1(18,44),
			in2                => s_in2(18,44),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(44)
		);
	s_in1(18,44)            <= s_out1(19,44);
	s_in2(18,44)            <= s_out2(19,45);
	s_locks_lower_in(18,44) <= s_locks_lower_out(19,44);

		normal_cell_18_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,45),
			fetch              => s_fetch(18,45),
			data_in            => s_data_in(18,45),
			data_out           => s_data_out(18,45),
			out1               => s_out1(18,45),
			out2               => s_out2(18,45),
			lock_lower_row_out => s_locks_lower_out(18,45),
			lock_lower_row_in  => s_locks_lower_in(18,45),
			in1                => s_in1(18,45),
			in2                => s_in2(18,45),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(45)
		);
	s_in1(18,45)            <= s_out1(19,45);
	s_in2(18,45)            <= s_out2(19,46);
	s_locks_lower_in(18,45) <= s_locks_lower_out(19,45);

		normal_cell_18_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,46),
			fetch              => s_fetch(18,46),
			data_in            => s_data_in(18,46),
			data_out           => s_data_out(18,46),
			out1               => s_out1(18,46),
			out2               => s_out2(18,46),
			lock_lower_row_out => s_locks_lower_out(18,46),
			lock_lower_row_in  => s_locks_lower_in(18,46),
			in1                => s_in1(18,46),
			in2                => s_in2(18,46),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(46)
		);
	s_in1(18,46)            <= s_out1(19,46);
	s_in2(18,46)            <= s_out2(19,47);
	s_locks_lower_in(18,46) <= s_locks_lower_out(19,46);

		normal_cell_18_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,47),
			fetch              => s_fetch(18,47),
			data_in            => s_data_in(18,47),
			data_out           => s_data_out(18,47),
			out1               => s_out1(18,47),
			out2               => s_out2(18,47),
			lock_lower_row_out => s_locks_lower_out(18,47),
			lock_lower_row_in  => s_locks_lower_in(18,47),
			in1                => s_in1(18,47),
			in2                => s_in2(18,47),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(47)
		);
	s_in1(18,47)            <= s_out1(19,47);
	s_in2(18,47)            <= s_out2(19,48);
	s_locks_lower_in(18,47) <= s_locks_lower_out(19,47);

		normal_cell_18_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,48),
			fetch              => s_fetch(18,48),
			data_in            => s_data_in(18,48),
			data_out           => s_data_out(18,48),
			out1               => s_out1(18,48),
			out2               => s_out2(18,48),
			lock_lower_row_out => s_locks_lower_out(18,48),
			lock_lower_row_in  => s_locks_lower_in(18,48),
			in1                => s_in1(18,48),
			in2                => s_in2(18,48),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(48)
		);
	s_in1(18,48)            <= s_out1(19,48);
	s_in2(18,48)            <= s_out2(19,49);
	s_locks_lower_in(18,48) <= s_locks_lower_out(19,48);

		normal_cell_18_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,49),
			fetch              => s_fetch(18,49),
			data_in            => s_data_in(18,49),
			data_out           => s_data_out(18,49),
			out1               => s_out1(18,49),
			out2               => s_out2(18,49),
			lock_lower_row_out => s_locks_lower_out(18,49),
			lock_lower_row_in  => s_locks_lower_in(18,49),
			in1                => s_in1(18,49),
			in2                => s_in2(18,49),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(49)
		);
	s_in1(18,49)            <= s_out1(19,49);
	s_in2(18,49)            <= s_out2(19,50);
	s_locks_lower_in(18,49) <= s_locks_lower_out(19,49);

		normal_cell_18_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,50),
			fetch              => s_fetch(18,50),
			data_in            => s_data_in(18,50),
			data_out           => s_data_out(18,50),
			out1               => s_out1(18,50),
			out2               => s_out2(18,50),
			lock_lower_row_out => s_locks_lower_out(18,50),
			lock_lower_row_in  => s_locks_lower_in(18,50),
			in1                => s_in1(18,50),
			in2                => s_in2(18,50),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(50)
		);
	s_in1(18,50)            <= s_out1(19,50);
	s_in2(18,50)            <= s_out2(19,51);
	s_locks_lower_in(18,50) <= s_locks_lower_out(19,50);

		normal_cell_18_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,51),
			fetch              => s_fetch(18,51),
			data_in            => s_data_in(18,51),
			data_out           => s_data_out(18,51),
			out1               => s_out1(18,51),
			out2               => s_out2(18,51),
			lock_lower_row_out => s_locks_lower_out(18,51),
			lock_lower_row_in  => s_locks_lower_in(18,51),
			in1                => s_in1(18,51),
			in2                => s_in2(18,51),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(51)
		);
	s_in1(18,51)            <= s_out1(19,51);
	s_in2(18,51)            <= s_out2(19,52);
	s_locks_lower_in(18,51) <= s_locks_lower_out(19,51);

		normal_cell_18_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,52),
			fetch              => s_fetch(18,52),
			data_in            => s_data_in(18,52),
			data_out           => s_data_out(18,52),
			out1               => s_out1(18,52),
			out2               => s_out2(18,52),
			lock_lower_row_out => s_locks_lower_out(18,52),
			lock_lower_row_in  => s_locks_lower_in(18,52),
			in1                => s_in1(18,52),
			in2                => s_in2(18,52),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(52)
		);
	s_in1(18,52)            <= s_out1(19,52);
	s_in2(18,52)            <= s_out2(19,53);
	s_locks_lower_in(18,52) <= s_locks_lower_out(19,52);

		normal_cell_18_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,53),
			fetch              => s_fetch(18,53),
			data_in            => s_data_in(18,53),
			data_out           => s_data_out(18,53),
			out1               => s_out1(18,53),
			out2               => s_out2(18,53),
			lock_lower_row_out => s_locks_lower_out(18,53),
			lock_lower_row_in  => s_locks_lower_in(18,53),
			in1                => s_in1(18,53),
			in2                => s_in2(18,53),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(53)
		);
	s_in1(18,53)            <= s_out1(19,53);
	s_in2(18,53)            <= s_out2(19,54);
	s_locks_lower_in(18,53) <= s_locks_lower_out(19,53);

		normal_cell_18_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,54),
			fetch              => s_fetch(18,54),
			data_in            => s_data_in(18,54),
			data_out           => s_data_out(18,54),
			out1               => s_out1(18,54),
			out2               => s_out2(18,54),
			lock_lower_row_out => s_locks_lower_out(18,54),
			lock_lower_row_in  => s_locks_lower_in(18,54),
			in1                => s_in1(18,54),
			in2                => s_in2(18,54),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(54)
		);
	s_in1(18,54)            <= s_out1(19,54);
	s_in2(18,54)            <= s_out2(19,55);
	s_locks_lower_in(18,54) <= s_locks_lower_out(19,54);

		normal_cell_18_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,55),
			fetch              => s_fetch(18,55),
			data_in            => s_data_in(18,55),
			data_out           => s_data_out(18,55),
			out1               => s_out1(18,55),
			out2               => s_out2(18,55),
			lock_lower_row_out => s_locks_lower_out(18,55),
			lock_lower_row_in  => s_locks_lower_in(18,55),
			in1                => s_in1(18,55),
			in2                => s_in2(18,55),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(55)
		);
	s_in1(18,55)            <= s_out1(19,55);
	s_in2(18,55)            <= s_out2(19,56);
	s_locks_lower_in(18,55) <= s_locks_lower_out(19,55);

		normal_cell_18_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,56),
			fetch              => s_fetch(18,56),
			data_in            => s_data_in(18,56),
			data_out           => s_data_out(18,56),
			out1               => s_out1(18,56),
			out2               => s_out2(18,56),
			lock_lower_row_out => s_locks_lower_out(18,56),
			lock_lower_row_in  => s_locks_lower_in(18,56),
			in1                => s_in1(18,56),
			in2                => s_in2(18,56),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(56)
		);
	s_in1(18,56)            <= s_out1(19,56);
	s_in2(18,56)            <= s_out2(19,57);
	s_locks_lower_in(18,56) <= s_locks_lower_out(19,56);

		normal_cell_18_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,57),
			fetch              => s_fetch(18,57),
			data_in            => s_data_in(18,57),
			data_out           => s_data_out(18,57),
			out1               => s_out1(18,57),
			out2               => s_out2(18,57),
			lock_lower_row_out => s_locks_lower_out(18,57),
			lock_lower_row_in  => s_locks_lower_in(18,57),
			in1                => s_in1(18,57),
			in2                => s_in2(18,57),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(57)
		);
	s_in1(18,57)            <= s_out1(19,57);
	s_in2(18,57)            <= s_out2(19,58);
	s_locks_lower_in(18,57) <= s_locks_lower_out(19,57);

		normal_cell_18_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,58),
			fetch              => s_fetch(18,58),
			data_in            => s_data_in(18,58),
			data_out           => s_data_out(18,58),
			out1               => s_out1(18,58),
			out2               => s_out2(18,58),
			lock_lower_row_out => s_locks_lower_out(18,58),
			lock_lower_row_in  => s_locks_lower_in(18,58),
			in1                => s_in1(18,58),
			in2                => s_in2(18,58),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(58)
		);
	s_in1(18,58)            <= s_out1(19,58);
	s_in2(18,58)            <= s_out2(19,59);
	s_locks_lower_in(18,58) <= s_locks_lower_out(19,58);

		normal_cell_18_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,59),
			fetch              => s_fetch(18,59),
			data_in            => s_data_in(18,59),
			data_out           => s_data_out(18,59),
			out1               => s_out1(18,59),
			out2               => s_out2(18,59),
			lock_lower_row_out => s_locks_lower_out(18,59),
			lock_lower_row_in  => s_locks_lower_in(18,59),
			in1                => s_in1(18,59),
			in2                => s_in2(18,59),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(59)
		);
	s_in1(18,59)            <= s_out1(19,59);
	s_in2(18,59)            <= s_out2(19,60);
	s_locks_lower_in(18,59) <= s_locks_lower_out(19,59);

		last_col_cell_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(18,60),
			fetch              => s_fetch(18,60),
			data_in            => s_data_in(18,60),
			data_out           => s_data_out(18,60),
			out1               => s_out1(18,60),
			out2               => s_out2(18,60),
			lock_lower_row_out => s_locks_lower_out(18,60),
			lock_lower_row_in  => s_locks_lower_in(18,60),
			in1                => s_in1(18,60),
			in2                => (others => '0'),
			lock_row           => s_locks(18),
			piv_found          => s_piv_found,
			row_data           => s_row_data(18),
			col_data           => s_col_data(60)
		);
	s_in1(18,60)            <= s_out1(19,60);
	s_locks_lower_in(18,60) <= s_locks_lower_out(19,60);

		normal_cell_19_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,1),
			fetch              => s_fetch(19,1),
			data_in            => s_data_in(19,1),
			data_out           => s_data_out(19,1),
			out1               => s_out1(19,1),
			out2               => s_out2(19,1),
			lock_lower_row_out => s_locks_lower_out(19,1),
			lock_lower_row_in  => s_locks_lower_in(19,1),
			in1                => s_in1(19,1),
			in2                => s_in2(19,1),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(1)
		);
	s_in1(19,1)            <= s_out1(20,1);
	s_in2(19,1)            <= s_out2(20,2);
	s_locks_lower_in(19,1) <= s_locks_lower_out(20,1);

		normal_cell_19_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,2),
			fetch              => s_fetch(19,2),
			data_in            => s_data_in(19,2),
			data_out           => s_data_out(19,2),
			out1               => s_out1(19,2),
			out2               => s_out2(19,2),
			lock_lower_row_out => s_locks_lower_out(19,2),
			lock_lower_row_in  => s_locks_lower_in(19,2),
			in1                => s_in1(19,2),
			in2                => s_in2(19,2),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(2)
		);
	s_in1(19,2)            <= s_out1(20,2);
	s_in2(19,2)            <= s_out2(20,3);
	s_locks_lower_in(19,2) <= s_locks_lower_out(20,2);

		normal_cell_19_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,3),
			fetch              => s_fetch(19,3),
			data_in            => s_data_in(19,3),
			data_out           => s_data_out(19,3),
			out1               => s_out1(19,3),
			out2               => s_out2(19,3),
			lock_lower_row_out => s_locks_lower_out(19,3),
			lock_lower_row_in  => s_locks_lower_in(19,3),
			in1                => s_in1(19,3),
			in2                => s_in2(19,3),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(3)
		);
	s_in1(19,3)            <= s_out1(20,3);
	s_in2(19,3)            <= s_out2(20,4);
	s_locks_lower_in(19,3) <= s_locks_lower_out(20,3);

		normal_cell_19_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,4),
			fetch              => s_fetch(19,4),
			data_in            => s_data_in(19,4),
			data_out           => s_data_out(19,4),
			out1               => s_out1(19,4),
			out2               => s_out2(19,4),
			lock_lower_row_out => s_locks_lower_out(19,4),
			lock_lower_row_in  => s_locks_lower_in(19,4),
			in1                => s_in1(19,4),
			in2                => s_in2(19,4),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(4)
		);
	s_in1(19,4)            <= s_out1(20,4);
	s_in2(19,4)            <= s_out2(20,5);
	s_locks_lower_in(19,4) <= s_locks_lower_out(20,4);

		normal_cell_19_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,5),
			fetch              => s_fetch(19,5),
			data_in            => s_data_in(19,5),
			data_out           => s_data_out(19,5),
			out1               => s_out1(19,5),
			out2               => s_out2(19,5),
			lock_lower_row_out => s_locks_lower_out(19,5),
			lock_lower_row_in  => s_locks_lower_in(19,5),
			in1                => s_in1(19,5),
			in2                => s_in2(19,5),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(5)
		);
	s_in1(19,5)            <= s_out1(20,5);
	s_in2(19,5)            <= s_out2(20,6);
	s_locks_lower_in(19,5) <= s_locks_lower_out(20,5);

		normal_cell_19_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,6),
			fetch              => s_fetch(19,6),
			data_in            => s_data_in(19,6),
			data_out           => s_data_out(19,6),
			out1               => s_out1(19,6),
			out2               => s_out2(19,6),
			lock_lower_row_out => s_locks_lower_out(19,6),
			lock_lower_row_in  => s_locks_lower_in(19,6),
			in1                => s_in1(19,6),
			in2                => s_in2(19,6),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(6)
		);
	s_in1(19,6)            <= s_out1(20,6);
	s_in2(19,6)            <= s_out2(20,7);
	s_locks_lower_in(19,6) <= s_locks_lower_out(20,6);

		normal_cell_19_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,7),
			fetch              => s_fetch(19,7),
			data_in            => s_data_in(19,7),
			data_out           => s_data_out(19,7),
			out1               => s_out1(19,7),
			out2               => s_out2(19,7),
			lock_lower_row_out => s_locks_lower_out(19,7),
			lock_lower_row_in  => s_locks_lower_in(19,7),
			in1                => s_in1(19,7),
			in2                => s_in2(19,7),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(7)
		);
	s_in1(19,7)            <= s_out1(20,7);
	s_in2(19,7)            <= s_out2(20,8);
	s_locks_lower_in(19,7) <= s_locks_lower_out(20,7);

		normal_cell_19_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,8),
			fetch              => s_fetch(19,8),
			data_in            => s_data_in(19,8),
			data_out           => s_data_out(19,8),
			out1               => s_out1(19,8),
			out2               => s_out2(19,8),
			lock_lower_row_out => s_locks_lower_out(19,8),
			lock_lower_row_in  => s_locks_lower_in(19,8),
			in1                => s_in1(19,8),
			in2                => s_in2(19,8),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(8)
		);
	s_in1(19,8)            <= s_out1(20,8);
	s_in2(19,8)            <= s_out2(20,9);
	s_locks_lower_in(19,8) <= s_locks_lower_out(20,8);

		normal_cell_19_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,9),
			fetch              => s_fetch(19,9),
			data_in            => s_data_in(19,9),
			data_out           => s_data_out(19,9),
			out1               => s_out1(19,9),
			out2               => s_out2(19,9),
			lock_lower_row_out => s_locks_lower_out(19,9),
			lock_lower_row_in  => s_locks_lower_in(19,9),
			in1                => s_in1(19,9),
			in2                => s_in2(19,9),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(9)
		);
	s_in1(19,9)            <= s_out1(20,9);
	s_in2(19,9)            <= s_out2(20,10);
	s_locks_lower_in(19,9) <= s_locks_lower_out(20,9);

		normal_cell_19_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,10),
			fetch              => s_fetch(19,10),
			data_in            => s_data_in(19,10),
			data_out           => s_data_out(19,10),
			out1               => s_out1(19,10),
			out2               => s_out2(19,10),
			lock_lower_row_out => s_locks_lower_out(19,10),
			lock_lower_row_in  => s_locks_lower_in(19,10),
			in1                => s_in1(19,10),
			in2                => s_in2(19,10),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(10)
		);
	s_in1(19,10)            <= s_out1(20,10);
	s_in2(19,10)            <= s_out2(20,11);
	s_locks_lower_in(19,10) <= s_locks_lower_out(20,10);

		normal_cell_19_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,11),
			fetch              => s_fetch(19,11),
			data_in            => s_data_in(19,11),
			data_out           => s_data_out(19,11),
			out1               => s_out1(19,11),
			out2               => s_out2(19,11),
			lock_lower_row_out => s_locks_lower_out(19,11),
			lock_lower_row_in  => s_locks_lower_in(19,11),
			in1                => s_in1(19,11),
			in2                => s_in2(19,11),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(11)
		);
	s_in1(19,11)            <= s_out1(20,11);
	s_in2(19,11)            <= s_out2(20,12);
	s_locks_lower_in(19,11) <= s_locks_lower_out(20,11);

		normal_cell_19_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,12),
			fetch              => s_fetch(19,12),
			data_in            => s_data_in(19,12),
			data_out           => s_data_out(19,12),
			out1               => s_out1(19,12),
			out2               => s_out2(19,12),
			lock_lower_row_out => s_locks_lower_out(19,12),
			lock_lower_row_in  => s_locks_lower_in(19,12),
			in1                => s_in1(19,12),
			in2                => s_in2(19,12),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(12)
		);
	s_in1(19,12)            <= s_out1(20,12);
	s_in2(19,12)            <= s_out2(20,13);
	s_locks_lower_in(19,12) <= s_locks_lower_out(20,12);

		normal_cell_19_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,13),
			fetch              => s_fetch(19,13),
			data_in            => s_data_in(19,13),
			data_out           => s_data_out(19,13),
			out1               => s_out1(19,13),
			out2               => s_out2(19,13),
			lock_lower_row_out => s_locks_lower_out(19,13),
			lock_lower_row_in  => s_locks_lower_in(19,13),
			in1                => s_in1(19,13),
			in2                => s_in2(19,13),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(13)
		);
	s_in1(19,13)            <= s_out1(20,13);
	s_in2(19,13)            <= s_out2(20,14);
	s_locks_lower_in(19,13) <= s_locks_lower_out(20,13);

		normal_cell_19_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,14),
			fetch              => s_fetch(19,14),
			data_in            => s_data_in(19,14),
			data_out           => s_data_out(19,14),
			out1               => s_out1(19,14),
			out2               => s_out2(19,14),
			lock_lower_row_out => s_locks_lower_out(19,14),
			lock_lower_row_in  => s_locks_lower_in(19,14),
			in1                => s_in1(19,14),
			in2                => s_in2(19,14),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(14)
		);
	s_in1(19,14)            <= s_out1(20,14);
	s_in2(19,14)            <= s_out2(20,15);
	s_locks_lower_in(19,14) <= s_locks_lower_out(20,14);

		normal_cell_19_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,15),
			fetch              => s_fetch(19,15),
			data_in            => s_data_in(19,15),
			data_out           => s_data_out(19,15),
			out1               => s_out1(19,15),
			out2               => s_out2(19,15),
			lock_lower_row_out => s_locks_lower_out(19,15),
			lock_lower_row_in  => s_locks_lower_in(19,15),
			in1                => s_in1(19,15),
			in2                => s_in2(19,15),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(15)
		);
	s_in1(19,15)            <= s_out1(20,15);
	s_in2(19,15)            <= s_out2(20,16);
	s_locks_lower_in(19,15) <= s_locks_lower_out(20,15);

		normal_cell_19_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,16),
			fetch              => s_fetch(19,16),
			data_in            => s_data_in(19,16),
			data_out           => s_data_out(19,16),
			out1               => s_out1(19,16),
			out2               => s_out2(19,16),
			lock_lower_row_out => s_locks_lower_out(19,16),
			lock_lower_row_in  => s_locks_lower_in(19,16),
			in1                => s_in1(19,16),
			in2                => s_in2(19,16),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(16)
		);
	s_in1(19,16)            <= s_out1(20,16);
	s_in2(19,16)            <= s_out2(20,17);
	s_locks_lower_in(19,16) <= s_locks_lower_out(20,16);

		normal_cell_19_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,17),
			fetch              => s_fetch(19,17),
			data_in            => s_data_in(19,17),
			data_out           => s_data_out(19,17),
			out1               => s_out1(19,17),
			out2               => s_out2(19,17),
			lock_lower_row_out => s_locks_lower_out(19,17),
			lock_lower_row_in  => s_locks_lower_in(19,17),
			in1                => s_in1(19,17),
			in2                => s_in2(19,17),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(17)
		);
	s_in1(19,17)            <= s_out1(20,17);
	s_in2(19,17)            <= s_out2(20,18);
	s_locks_lower_in(19,17) <= s_locks_lower_out(20,17);

		normal_cell_19_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,18),
			fetch              => s_fetch(19,18),
			data_in            => s_data_in(19,18),
			data_out           => s_data_out(19,18),
			out1               => s_out1(19,18),
			out2               => s_out2(19,18),
			lock_lower_row_out => s_locks_lower_out(19,18),
			lock_lower_row_in  => s_locks_lower_in(19,18),
			in1                => s_in1(19,18),
			in2                => s_in2(19,18),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(18)
		);
	s_in1(19,18)            <= s_out1(20,18);
	s_in2(19,18)            <= s_out2(20,19);
	s_locks_lower_in(19,18) <= s_locks_lower_out(20,18);

		normal_cell_19_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,19),
			fetch              => s_fetch(19,19),
			data_in            => s_data_in(19,19),
			data_out           => s_data_out(19,19),
			out1               => s_out1(19,19),
			out2               => s_out2(19,19),
			lock_lower_row_out => s_locks_lower_out(19,19),
			lock_lower_row_in  => s_locks_lower_in(19,19),
			in1                => s_in1(19,19),
			in2                => s_in2(19,19),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(19)
		);
	s_in1(19,19)            <= s_out1(20,19);
	s_in2(19,19)            <= s_out2(20,20);
	s_locks_lower_in(19,19) <= s_locks_lower_out(20,19);

		normal_cell_19_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,20),
			fetch              => s_fetch(19,20),
			data_in            => s_data_in(19,20),
			data_out           => s_data_out(19,20),
			out1               => s_out1(19,20),
			out2               => s_out2(19,20),
			lock_lower_row_out => s_locks_lower_out(19,20),
			lock_lower_row_in  => s_locks_lower_in(19,20),
			in1                => s_in1(19,20),
			in2                => s_in2(19,20),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(20)
		);
	s_in1(19,20)            <= s_out1(20,20);
	s_in2(19,20)            <= s_out2(20,21);
	s_locks_lower_in(19,20) <= s_locks_lower_out(20,20);

		normal_cell_19_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,21),
			fetch              => s_fetch(19,21),
			data_in            => s_data_in(19,21),
			data_out           => s_data_out(19,21),
			out1               => s_out1(19,21),
			out2               => s_out2(19,21),
			lock_lower_row_out => s_locks_lower_out(19,21),
			lock_lower_row_in  => s_locks_lower_in(19,21),
			in1                => s_in1(19,21),
			in2                => s_in2(19,21),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(21)
		);
	s_in1(19,21)            <= s_out1(20,21);
	s_in2(19,21)            <= s_out2(20,22);
	s_locks_lower_in(19,21) <= s_locks_lower_out(20,21);

		normal_cell_19_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,22),
			fetch              => s_fetch(19,22),
			data_in            => s_data_in(19,22),
			data_out           => s_data_out(19,22),
			out1               => s_out1(19,22),
			out2               => s_out2(19,22),
			lock_lower_row_out => s_locks_lower_out(19,22),
			lock_lower_row_in  => s_locks_lower_in(19,22),
			in1                => s_in1(19,22),
			in2                => s_in2(19,22),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(22)
		);
	s_in1(19,22)            <= s_out1(20,22);
	s_in2(19,22)            <= s_out2(20,23);
	s_locks_lower_in(19,22) <= s_locks_lower_out(20,22);

		normal_cell_19_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,23),
			fetch              => s_fetch(19,23),
			data_in            => s_data_in(19,23),
			data_out           => s_data_out(19,23),
			out1               => s_out1(19,23),
			out2               => s_out2(19,23),
			lock_lower_row_out => s_locks_lower_out(19,23),
			lock_lower_row_in  => s_locks_lower_in(19,23),
			in1                => s_in1(19,23),
			in2                => s_in2(19,23),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(23)
		);
	s_in1(19,23)            <= s_out1(20,23);
	s_in2(19,23)            <= s_out2(20,24);
	s_locks_lower_in(19,23) <= s_locks_lower_out(20,23);

		normal_cell_19_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,24),
			fetch              => s_fetch(19,24),
			data_in            => s_data_in(19,24),
			data_out           => s_data_out(19,24),
			out1               => s_out1(19,24),
			out2               => s_out2(19,24),
			lock_lower_row_out => s_locks_lower_out(19,24),
			lock_lower_row_in  => s_locks_lower_in(19,24),
			in1                => s_in1(19,24),
			in2                => s_in2(19,24),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(24)
		);
	s_in1(19,24)            <= s_out1(20,24);
	s_in2(19,24)            <= s_out2(20,25);
	s_locks_lower_in(19,24) <= s_locks_lower_out(20,24);

		normal_cell_19_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,25),
			fetch              => s_fetch(19,25),
			data_in            => s_data_in(19,25),
			data_out           => s_data_out(19,25),
			out1               => s_out1(19,25),
			out2               => s_out2(19,25),
			lock_lower_row_out => s_locks_lower_out(19,25),
			lock_lower_row_in  => s_locks_lower_in(19,25),
			in1                => s_in1(19,25),
			in2                => s_in2(19,25),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(25)
		);
	s_in1(19,25)            <= s_out1(20,25);
	s_in2(19,25)            <= s_out2(20,26);
	s_locks_lower_in(19,25) <= s_locks_lower_out(20,25);

		normal_cell_19_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,26),
			fetch              => s_fetch(19,26),
			data_in            => s_data_in(19,26),
			data_out           => s_data_out(19,26),
			out1               => s_out1(19,26),
			out2               => s_out2(19,26),
			lock_lower_row_out => s_locks_lower_out(19,26),
			lock_lower_row_in  => s_locks_lower_in(19,26),
			in1                => s_in1(19,26),
			in2                => s_in2(19,26),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(26)
		);
	s_in1(19,26)            <= s_out1(20,26);
	s_in2(19,26)            <= s_out2(20,27);
	s_locks_lower_in(19,26) <= s_locks_lower_out(20,26);

		normal_cell_19_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,27),
			fetch              => s_fetch(19,27),
			data_in            => s_data_in(19,27),
			data_out           => s_data_out(19,27),
			out1               => s_out1(19,27),
			out2               => s_out2(19,27),
			lock_lower_row_out => s_locks_lower_out(19,27),
			lock_lower_row_in  => s_locks_lower_in(19,27),
			in1                => s_in1(19,27),
			in2                => s_in2(19,27),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(27)
		);
	s_in1(19,27)            <= s_out1(20,27);
	s_in2(19,27)            <= s_out2(20,28);
	s_locks_lower_in(19,27) <= s_locks_lower_out(20,27);

		normal_cell_19_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,28),
			fetch              => s_fetch(19,28),
			data_in            => s_data_in(19,28),
			data_out           => s_data_out(19,28),
			out1               => s_out1(19,28),
			out2               => s_out2(19,28),
			lock_lower_row_out => s_locks_lower_out(19,28),
			lock_lower_row_in  => s_locks_lower_in(19,28),
			in1                => s_in1(19,28),
			in2                => s_in2(19,28),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(28)
		);
	s_in1(19,28)            <= s_out1(20,28);
	s_in2(19,28)            <= s_out2(20,29);
	s_locks_lower_in(19,28) <= s_locks_lower_out(20,28);

		normal_cell_19_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,29),
			fetch              => s_fetch(19,29),
			data_in            => s_data_in(19,29),
			data_out           => s_data_out(19,29),
			out1               => s_out1(19,29),
			out2               => s_out2(19,29),
			lock_lower_row_out => s_locks_lower_out(19,29),
			lock_lower_row_in  => s_locks_lower_in(19,29),
			in1                => s_in1(19,29),
			in2                => s_in2(19,29),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(29)
		);
	s_in1(19,29)            <= s_out1(20,29);
	s_in2(19,29)            <= s_out2(20,30);
	s_locks_lower_in(19,29) <= s_locks_lower_out(20,29);

		normal_cell_19_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,30),
			fetch              => s_fetch(19,30),
			data_in            => s_data_in(19,30),
			data_out           => s_data_out(19,30),
			out1               => s_out1(19,30),
			out2               => s_out2(19,30),
			lock_lower_row_out => s_locks_lower_out(19,30),
			lock_lower_row_in  => s_locks_lower_in(19,30),
			in1                => s_in1(19,30),
			in2                => s_in2(19,30),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(30)
		);
	s_in1(19,30)            <= s_out1(20,30);
	s_in2(19,30)            <= s_out2(20,31);
	s_locks_lower_in(19,30) <= s_locks_lower_out(20,30);

		normal_cell_19_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,31),
			fetch              => s_fetch(19,31),
			data_in            => s_data_in(19,31),
			data_out           => s_data_out(19,31),
			out1               => s_out1(19,31),
			out2               => s_out2(19,31),
			lock_lower_row_out => s_locks_lower_out(19,31),
			lock_lower_row_in  => s_locks_lower_in(19,31),
			in1                => s_in1(19,31),
			in2                => s_in2(19,31),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(31)
		);
	s_in1(19,31)            <= s_out1(20,31);
	s_in2(19,31)            <= s_out2(20,32);
	s_locks_lower_in(19,31) <= s_locks_lower_out(20,31);

		normal_cell_19_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,32),
			fetch              => s_fetch(19,32),
			data_in            => s_data_in(19,32),
			data_out           => s_data_out(19,32),
			out1               => s_out1(19,32),
			out2               => s_out2(19,32),
			lock_lower_row_out => s_locks_lower_out(19,32),
			lock_lower_row_in  => s_locks_lower_in(19,32),
			in1                => s_in1(19,32),
			in2                => s_in2(19,32),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(32)
		);
	s_in1(19,32)            <= s_out1(20,32);
	s_in2(19,32)            <= s_out2(20,33);
	s_locks_lower_in(19,32) <= s_locks_lower_out(20,32);

		normal_cell_19_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,33),
			fetch              => s_fetch(19,33),
			data_in            => s_data_in(19,33),
			data_out           => s_data_out(19,33),
			out1               => s_out1(19,33),
			out2               => s_out2(19,33),
			lock_lower_row_out => s_locks_lower_out(19,33),
			lock_lower_row_in  => s_locks_lower_in(19,33),
			in1                => s_in1(19,33),
			in2                => s_in2(19,33),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(33)
		);
	s_in1(19,33)            <= s_out1(20,33);
	s_in2(19,33)            <= s_out2(20,34);
	s_locks_lower_in(19,33) <= s_locks_lower_out(20,33);

		normal_cell_19_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,34),
			fetch              => s_fetch(19,34),
			data_in            => s_data_in(19,34),
			data_out           => s_data_out(19,34),
			out1               => s_out1(19,34),
			out2               => s_out2(19,34),
			lock_lower_row_out => s_locks_lower_out(19,34),
			lock_lower_row_in  => s_locks_lower_in(19,34),
			in1                => s_in1(19,34),
			in2                => s_in2(19,34),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(34)
		);
	s_in1(19,34)            <= s_out1(20,34);
	s_in2(19,34)            <= s_out2(20,35);
	s_locks_lower_in(19,34) <= s_locks_lower_out(20,34);

		normal_cell_19_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,35),
			fetch              => s_fetch(19,35),
			data_in            => s_data_in(19,35),
			data_out           => s_data_out(19,35),
			out1               => s_out1(19,35),
			out2               => s_out2(19,35),
			lock_lower_row_out => s_locks_lower_out(19,35),
			lock_lower_row_in  => s_locks_lower_in(19,35),
			in1                => s_in1(19,35),
			in2                => s_in2(19,35),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(35)
		);
	s_in1(19,35)            <= s_out1(20,35);
	s_in2(19,35)            <= s_out2(20,36);
	s_locks_lower_in(19,35) <= s_locks_lower_out(20,35);

		normal_cell_19_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,36),
			fetch              => s_fetch(19,36),
			data_in            => s_data_in(19,36),
			data_out           => s_data_out(19,36),
			out1               => s_out1(19,36),
			out2               => s_out2(19,36),
			lock_lower_row_out => s_locks_lower_out(19,36),
			lock_lower_row_in  => s_locks_lower_in(19,36),
			in1                => s_in1(19,36),
			in2                => s_in2(19,36),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(36)
		);
	s_in1(19,36)            <= s_out1(20,36);
	s_in2(19,36)            <= s_out2(20,37);
	s_locks_lower_in(19,36) <= s_locks_lower_out(20,36);

		normal_cell_19_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,37),
			fetch              => s_fetch(19,37),
			data_in            => s_data_in(19,37),
			data_out           => s_data_out(19,37),
			out1               => s_out1(19,37),
			out2               => s_out2(19,37),
			lock_lower_row_out => s_locks_lower_out(19,37),
			lock_lower_row_in  => s_locks_lower_in(19,37),
			in1                => s_in1(19,37),
			in2                => s_in2(19,37),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(37)
		);
	s_in1(19,37)            <= s_out1(20,37);
	s_in2(19,37)            <= s_out2(20,38);
	s_locks_lower_in(19,37) <= s_locks_lower_out(20,37);

		normal_cell_19_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,38),
			fetch              => s_fetch(19,38),
			data_in            => s_data_in(19,38),
			data_out           => s_data_out(19,38),
			out1               => s_out1(19,38),
			out2               => s_out2(19,38),
			lock_lower_row_out => s_locks_lower_out(19,38),
			lock_lower_row_in  => s_locks_lower_in(19,38),
			in1                => s_in1(19,38),
			in2                => s_in2(19,38),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(38)
		);
	s_in1(19,38)            <= s_out1(20,38);
	s_in2(19,38)            <= s_out2(20,39);
	s_locks_lower_in(19,38) <= s_locks_lower_out(20,38);

		normal_cell_19_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,39),
			fetch              => s_fetch(19,39),
			data_in            => s_data_in(19,39),
			data_out           => s_data_out(19,39),
			out1               => s_out1(19,39),
			out2               => s_out2(19,39),
			lock_lower_row_out => s_locks_lower_out(19,39),
			lock_lower_row_in  => s_locks_lower_in(19,39),
			in1                => s_in1(19,39),
			in2                => s_in2(19,39),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(39)
		);
	s_in1(19,39)            <= s_out1(20,39);
	s_in2(19,39)            <= s_out2(20,40);
	s_locks_lower_in(19,39) <= s_locks_lower_out(20,39);

		normal_cell_19_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,40),
			fetch              => s_fetch(19,40),
			data_in            => s_data_in(19,40),
			data_out           => s_data_out(19,40),
			out1               => s_out1(19,40),
			out2               => s_out2(19,40),
			lock_lower_row_out => s_locks_lower_out(19,40),
			lock_lower_row_in  => s_locks_lower_in(19,40),
			in1                => s_in1(19,40),
			in2                => s_in2(19,40),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(40)
		);
	s_in1(19,40)            <= s_out1(20,40);
	s_in2(19,40)            <= s_out2(20,41);
	s_locks_lower_in(19,40) <= s_locks_lower_out(20,40);

		normal_cell_19_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,41),
			fetch              => s_fetch(19,41),
			data_in            => s_data_in(19,41),
			data_out           => s_data_out(19,41),
			out1               => s_out1(19,41),
			out2               => s_out2(19,41),
			lock_lower_row_out => s_locks_lower_out(19,41),
			lock_lower_row_in  => s_locks_lower_in(19,41),
			in1                => s_in1(19,41),
			in2                => s_in2(19,41),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(41)
		);
	s_in1(19,41)            <= s_out1(20,41);
	s_in2(19,41)            <= s_out2(20,42);
	s_locks_lower_in(19,41) <= s_locks_lower_out(20,41);

		normal_cell_19_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,42),
			fetch              => s_fetch(19,42),
			data_in            => s_data_in(19,42),
			data_out           => s_data_out(19,42),
			out1               => s_out1(19,42),
			out2               => s_out2(19,42),
			lock_lower_row_out => s_locks_lower_out(19,42),
			lock_lower_row_in  => s_locks_lower_in(19,42),
			in1                => s_in1(19,42),
			in2                => s_in2(19,42),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(42)
		);
	s_in1(19,42)            <= s_out1(20,42);
	s_in2(19,42)            <= s_out2(20,43);
	s_locks_lower_in(19,42) <= s_locks_lower_out(20,42);

		normal_cell_19_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,43),
			fetch              => s_fetch(19,43),
			data_in            => s_data_in(19,43),
			data_out           => s_data_out(19,43),
			out1               => s_out1(19,43),
			out2               => s_out2(19,43),
			lock_lower_row_out => s_locks_lower_out(19,43),
			lock_lower_row_in  => s_locks_lower_in(19,43),
			in1                => s_in1(19,43),
			in2                => s_in2(19,43),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(43)
		);
	s_in1(19,43)            <= s_out1(20,43);
	s_in2(19,43)            <= s_out2(20,44);
	s_locks_lower_in(19,43) <= s_locks_lower_out(20,43);

		normal_cell_19_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,44),
			fetch              => s_fetch(19,44),
			data_in            => s_data_in(19,44),
			data_out           => s_data_out(19,44),
			out1               => s_out1(19,44),
			out2               => s_out2(19,44),
			lock_lower_row_out => s_locks_lower_out(19,44),
			lock_lower_row_in  => s_locks_lower_in(19,44),
			in1                => s_in1(19,44),
			in2                => s_in2(19,44),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(44)
		);
	s_in1(19,44)            <= s_out1(20,44);
	s_in2(19,44)            <= s_out2(20,45);
	s_locks_lower_in(19,44) <= s_locks_lower_out(20,44);

		normal_cell_19_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,45),
			fetch              => s_fetch(19,45),
			data_in            => s_data_in(19,45),
			data_out           => s_data_out(19,45),
			out1               => s_out1(19,45),
			out2               => s_out2(19,45),
			lock_lower_row_out => s_locks_lower_out(19,45),
			lock_lower_row_in  => s_locks_lower_in(19,45),
			in1                => s_in1(19,45),
			in2                => s_in2(19,45),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(45)
		);
	s_in1(19,45)            <= s_out1(20,45);
	s_in2(19,45)            <= s_out2(20,46);
	s_locks_lower_in(19,45) <= s_locks_lower_out(20,45);

		normal_cell_19_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,46),
			fetch              => s_fetch(19,46),
			data_in            => s_data_in(19,46),
			data_out           => s_data_out(19,46),
			out1               => s_out1(19,46),
			out2               => s_out2(19,46),
			lock_lower_row_out => s_locks_lower_out(19,46),
			lock_lower_row_in  => s_locks_lower_in(19,46),
			in1                => s_in1(19,46),
			in2                => s_in2(19,46),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(46)
		);
	s_in1(19,46)            <= s_out1(20,46);
	s_in2(19,46)            <= s_out2(20,47);
	s_locks_lower_in(19,46) <= s_locks_lower_out(20,46);

		normal_cell_19_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,47),
			fetch              => s_fetch(19,47),
			data_in            => s_data_in(19,47),
			data_out           => s_data_out(19,47),
			out1               => s_out1(19,47),
			out2               => s_out2(19,47),
			lock_lower_row_out => s_locks_lower_out(19,47),
			lock_lower_row_in  => s_locks_lower_in(19,47),
			in1                => s_in1(19,47),
			in2                => s_in2(19,47),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(47)
		);
	s_in1(19,47)            <= s_out1(20,47);
	s_in2(19,47)            <= s_out2(20,48);
	s_locks_lower_in(19,47) <= s_locks_lower_out(20,47);

		normal_cell_19_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,48),
			fetch              => s_fetch(19,48),
			data_in            => s_data_in(19,48),
			data_out           => s_data_out(19,48),
			out1               => s_out1(19,48),
			out2               => s_out2(19,48),
			lock_lower_row_out => s_locks_lower_out(19,48),
			lock_lower_row_in  => s_locks_lower_in(19,48),
			in1                => s_in1(19,48),
			in2                => s_in2(19,48),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(48)
		);
	s_in1(19,48)            <= s_out1(20,48);
	s_in2(19,48)            <= s_out2(20,49);
	s_locks_lower_in(19,48) <= s_locks_lower_out(20,48);

		normal_cell_19_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,49),
			fetch              => s_fetch(19,49),
			data_in            => s_data_in(19,49),
			data_out           => s_data_out(19,49),
			out1               => s_out1(19,49),
			out2               => s_out2(19,49),
			lock_lower_row_out => s_locks_lower_out(19,49),
			lock_lower_row_in  => s_locks_lower_in(19,49),
			in1                => s_in1(19,49),
			in2                => s_in2(19,49),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(49)
		);
	s_in1(19,49)            <= s_out1(20,49);
	s_in2(19,49)            <= s_out2(20,50);
	s_locks_lower_in(19,49) <= s_locks_lower_out(20,49);

		normal_cell_19_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,50),
			fetch              => s_fetch(19,50),
			data_in            => s_data_in(19,50),
			data_out           => s_data_out(19,50),
			out1               => s_out1(19,50),
			out2               => s_out2(19,50),
			lock_lower_row_out => s_locks_lower_out(19,50),
			lock_lower_row_in  => s_locks_lower_in(19,50),
			in1                => s_in1(19,50),
			in2                => s_in2(19,50),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(50)
		);
	s_in1(19,50)            <= s_out1(20,50);
	s_in2(19,50)            <= s_out2(20,51);
	s_locks_lower_in(19,50) <= s_locks_lower_out(20,50);

		normal_cell_19_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,51),
			fetch              => s_fetch(19,51),
			data_in            => s_data_in(19,51),
			data_out           => s_data_out(19,51),
			out1               => s_out1(19,51),
			out2               => s_out2(19,51),
			lock_lower_row_out => s_locks_lower_out(19,51),
			lock_lower_row_in  => s_locks_lower_in(19,51),
			in1                => s_in1(19,51),
			in2                => s_in2(19,51),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(51)
		);
	s_in1(19,51)            <= s_out1(20,51);
	s_in2(19,51)            <= s_out2(20,52);
	s_locks_lower_in(19,51) <= s_locks_lower_out(20,51);

		normal_cell_19_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,52),
			fetch              => s_fetch(19,52),
			data_in            => s_data_in(19,52),
			data_out           => s_data_out(19,52),
			out1               => s_out1(19,52),
			out2               => s_out2(19,52),
			lock_lower_row_out => s_locks_lower_out(19,52),
			lock_lower_row_in  => s_locks_lower_in(19,52),
			in1                => s_in1(19,52),
			in2                => s_in2(19,52),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(52)
		);
	s_in1(19,52)            <= s_out1(20,52);
	s_in2(19,52)            <= s_out2(20,53);
	s_locks_lower_in(19,52) <= s_locks_lower_out(20,52);

		normal_cell_19_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,53),
			fetch              => s_fetch(19,53),
			data_in            => s_data_in(19,53),
			data_out           => s_data_out(19,53),
			out1               => s_out1(19,53),
			out2               => s_out2(19,53),
			lock_lower_row_out => s_locks_lower_out(19,53),
			lock_lower_row_in  => s_locks_lower_in(19,53),
			in1                => s_in1(19,53),
			in2                => s_in2(19,53),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(53)
		);
	s_in1(19,53)            <= s_out1(20,53);
	s_in2(19,53)            <= s_out2(20,54);
	s_locks_lower_in(19,53) <= s_locks_lower_out(20,53);

		normal_cell_19_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,54),
			fetch              => s_fetch(19,54),
			data_in            => s_data_in(19,54),
			data_out           => s_data_out(19,54),
			out1               => s_out1(19,54),
			out2               => s_out2(19,54),
			lock_lower_row_out => s_locks_lower_out(19,54),
			lock_lower_row_in  => s_locks_lower_in(19,54),
			in1                => s_in1(19,54),
			in2                => s_in2(19,54),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(54)
		);
	s_in1(19,54)            <= s_out1(20,54);
	s_in2(19,54)            <= s_out2(20,55);
	s_locks_lower_in(19,54) <= s_locks_lower_out(20,54);

		normal_cell_19_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,55),
			fetch              => s_fetch(19,55),
			data_in            => s_data_in(19,55),
			data_out           => s_data_out(19,55),
			out1               => s_out1(19,55),
			out2               => s_out2(19,55),
			lock_lower_row_out => s_locks_lower_out(19,55),
			lock_lower_row_in  => s_locks_lower_in(19,55),
			in1                => s_in1(19,55),
			in2                => s_in2(19,55),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(55)
		);
	s_in1(19,55)            <= s_out1(20,55);
	s_in2(19,55)            <= s_out2(20,56);
	s_locks_lower_in(19,55) <= s_locks_lower_out(20,55);

		normal_cell_19_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,56),
			fetch              => s_fetch(19,56),
			data_in            => s_data_in(19,56),
			data_out           => s_data_out(19,56),
			out1               => s_out1(19,56),
			out2               => s_out2(19,56),
			lock_lower_row_out => s_locks_lower_out(19,56),
			lock_lower_row_in  => s_locks_lower_in(19,56),
			in1                => s_in1(19,56),
			in2                => s_in2(19,56),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(56)
		);
	s_in1(19,56)            <= s_out1(20,56);
	s_in2(19,56)            <= s_out2(20,57);
	s_locks_lower_in(19,56) <= s_locks_lower_out(20,56);

		normal_cell_19_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,57),
			fetch              => s_fetch(19,57),
			data_in            => s_data_in(19,57),
			data_out           => s_data_out(19,57),
			out1               => s_out1(19,57),
			out2               => s_out2(19,57),
			lock_lower_row_out => s_locks_lower_out(19,57),
			lock_lower_row_in  => s_locks_lower_in(19,57),
			in1                => s_in1(19,57),
			in2                => s_in2(19,57),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(57)
		);
	s_in1(19,57)            <= s_out1(20,57);
	s_in2(19,57)            <= s_out2(20,58);
	s_locks_lower_in(19,57) <= s_locks_lower_out(20,57);

		normal_cell_19_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,58),
			fetch              => s_fetch(19,58),
			data_in            => s_data_in(19,58),
			data_out           => s_data_out(19,58),
			out1               => s_out1(19,58),
			out2               => s_out2(19,58),
			lock_lower_row_out => s_locks_lower_out(19,58),
			lock_lower_row_in  => s_locks_lower_in(19,58),
			in1                => s_in1(19,58),
			in2                => s_in2(19,58),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(58)
		);
	s_in1(19,58)            <= s_out1(20,58);
	s_in2(19,58)            <= s_out2(20,59);
	s_locks_lower_in(19,58) <= s_locks_lower_out(20,58);

		normal_cell_19_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,59),
			fetch              => s_fetch(19,59),
			data_in            => s_data_in(19,59),
			data_out           => s_data_out(19,59),
			out1               => s_out1(19,59),
			out2               => s_out2(19,59),
			lock_lower_row_out => s_locks_lower_out(19,59),
			lock_lower_row_in  => s_locks_lower_in(19,59),
			in1                => s_in1(19,59),
			in2                => s_in2(19,59),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(59)
		);
	s_in1(19,59)            <= s_out1(20,59);
	s_in2(19,59)            <= s_out2(20,60);
	s_locks_lower_in(19,59) <= s_locks_lower_out(20,59);

		last_col_cell_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(19,60),
			fetch              => s_fetch(19,60),
			data_in            => s_data_in(19,60),
			data_out           => s_data_out(19,60),
			out1               => s_out1(19,60),
			out2               => s_out2(19,60),
			lock_lower_row_out => s_locks_lower_out(19,60),
			lock_lower_row_in  => s_locks_lower_in(19,60),
			in1                => s_in1(19,60),
			in2                => (others => '0'),
			lock_row           => s_locks(19),
			piv_found          => s_piv_found,
			row_data           => s_row_data(19),
			col_data           => s_col_data(60)
		);
	s_in1(19,60)            <= s_out1(20,60);
	s_locks_lower_in(19,60) <= s_locks_lower_out(20,60);

		normal_cell_20_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,1),
			fetch              => s_fetch(20,1),
			data_in            => s_data_in(20,1),
			data_out           => s_data_out(20,1),
			out1               => s_out1(20,1),
			out2               => s_out2(20,1),
			lock_lower_row_out => s_locks_lower_out(20,1),
			lock_lower_row_in  => s_locks_lower_in(20,1),
			in1                => s_in1(20,1),
			in2                => s_in2(20,1),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(1)
		);
	s_in1(20,1)            <= s_out1(21,1);
	s_in2(20,1)            <= s_out2(21,2);
	s_locks_lower_in(20,1) <= s_locks_lower_out(21,1);

		normal_cell_20_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,2),
			fetch              => s_fetch(20,2),
			data_in            => s_data_in(20,2),
			data_out           => s_data_out(20,2),
			out1               => s_out1(20,2),
			out2               => s_out2(20,2),
			lock_lower_row_out => s_locks_lower_out(20,2),
			lock_lower_row_in  => s_locks_lower_in(20,2),
			in1                => s_in1(20,2),
			in2                => s_in2(20,2),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(2)
		);
	s_in1(20,2)            <= s_out1(21,2);
	s_in2(20,2)            <= s_out2(21,3);
	s_locks_lower_in(20,2) <= s_locks_lower_out(21,2);

		normal_cell_20_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,3),
			fetch              => s_fetch(20,3),
			data_in            => s_data_in(20,3),
			data_out           => s_data_out(20,3),
			out1               => s_out1(20,3),
			out2               => s_out2(20,3),
			lock_lower_row_out => s_locks_lower_out(20,3),
			lock_lower_row_in  => s_locks_lower_in(20,3),
			in1                => s_in1(20,3),
			in2                => s_in2(20,3),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(3)
		);
	s_in1(20,3)            <= s_out1(21,3);
	s_in2(20,3)            <= s_out2(21,4);
	s_locks_lower_in(20,3) <= s_locks_lower_out(21,3);

		normal_cell_20_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,4),
			fetch              => s_fetch(20,4),
			data_in            => s_data_in(20,4),
			data_out           => s_data_out(20,4),
			out1               => s_out1(20,4),
			out2               => s_out2(20,4),
			lock_lower_row_out => s_locks_lower_out(20,4),
			lock_lower_row_in  => s_locks_lower_in(20,4),
			in1                => s_in1(20,4),
			in2                => s_in2(20,4),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(4)
		);
	s_in1(20,4)            <= s_out1(21,4);
	s_in2(20,4)            <= s_out2(21,5);
	s_locks_lower_in(20,4) <= s_locks_lower_out(21,4);

		normal_cell_20_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,5),
			fetch              => s_fetch(20,5),
			data_in            => s_data_in(20,5),
			data_out           => s_data_out(20,5),
			out1               => s_out1(20,5),
			out2               => s_out2(20,5),
			lock_lower_row_out => s_locks_lower_out(20,5),
			lock_lower_row_in  => s_locks_lower_in(20,5),
			in1                => s_in1(20,5),
			in2                => s_in2(20,5),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(5)
		);
	s_in1(20,5)            <= s_out1(21,5);
	s_in2(20,5)            <= s_out2(21,6);
	s_locks_lower_in(20,5) <= s_locks_lower_out(21,5);

		normal_cell_20_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,6),
			fetch              => s_fetch(20,6),
			data_in            => s_data_in(20,6),
			data_out           => s_data_out(20,6),
			out1               => s_out1(20,6),
			out2               => s_out2(20,6),
			lock_lower_row_out => s_locks_lower_out(20,6),
			lock_lower_row_in  => s_locks_lower_in(20,6),
			in1                => s_in1(20,6),
			in2                => s_in2(20,6),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(6)
		);
	s_in1(20,6)            <= s_out1(21,6);
	s_in2(20,6)            <= s_out2(21,7);
	s_locks_lower_in(20,6) <= s_locks_lower_out(21,6);

		normal_cell_20_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,7),
			fetch              => s_fetch(20,7),
			data_in            => s_data_in(20,7),
			data_out           => s_data_out(20,7),
			out1               => s_out1(20,7),
			out2               => s_out2(20,7),
			lock_lower_row_out => s_locks_lower_out(20,7),
			lock_lower_row_in  => s_locks_lower_in(20,7),
			in1                => s_in1(20,7),
			in2                => s_in2(20,7),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(7)
		);
	s_in1(20,7)            <= s_out1(21,7);
	s_in2(20,7)            <= s_out2(21,8);
	s_locks_lower_in(20,7) <= s_locks_lower_out(21,7);

		normal_cell_20_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,8),
			fetch              => s_fetch(20,8),
			data_in            => s_data_in(20,8),
			data_out           => s_data_out(20,8),
			out1               => s_out1(20,8),
			out2               => s_out2(20,8),
			lock_lower_row_out => s_locks_lower_out(20,8),
			lock_lower_row_in  => s_locks_lower_in(20,8),
			in1                => s_in1(20,8),
			in2                => s_in2(20,8),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(8)
		);
	s_in1(20,8)            <= s_out1(21,8);
	s_in2(20,8)            <= s_out2(21,9);
	s_locks_lower_in(20,8) <= s_locks_lower_out(21,8);

		normal_cell_20_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,9),
			fetch              => s_fetch(20,9),
			data_in            => s_data_in(20,9),
			data_out           => s_data_out(20,9),
			out1               => s_out1(20,9),
			out2               => s_out2(20,9),
			lock_lower_row_out => s_locks_lower_out(20,9),
			lock_lower_row_in  => s_locks_lower_in(20,9),
			in1                => s_in1(20,9),
			in2                => s_in2(20,9),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(9)
		);
	s_in1(20,9)            <= s_out1(21,9);
	s_in2(20,9)            <= s_out2(21,10);
	s_locks_lower_in(20,9) <= s_locks_lower_out(21,9);

		normal_cell_20_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,10),
			fetch              => s_fetch(20,10),
			data_in            => s_data_in(20,10),
			data_out           => s_data_out(20,10),
			out1               => s_out1(20,10),
			out2               => s_out2(20,10),
			lock_lower_row_out => s_locks_lower_out(20,10),
			lock_lower_row_in  => s_locks_lower_in(20,10),
			in1                => s_in1(20,10),
			in2                => s_in2(20,10),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(10)
		);
	s_in1(20,10)            <= s_out1(21,10);
	s_in2(20,10)            <= s_out2(21,11);
	s_locks_lower_in(20,10) <= s_locks_lower_out(21,10);

		normal_cell_20_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,11),
			fetch              => s_fetch(20,11),
			data_in            => s_data_in(20,11),
			data_out           => s_data_out(20,11),
			out1               => s_out1(20,11),
			out2               => s_out2(20,11),
			lock_lower_row_out => s_locks_lower_out(20,11),
			lock_lower_row_in  => s_locks_lower_in(20,11),
			in1                => s_in1(20,11),
			in2                => s_in2(20,11),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(11)
		);
	s_in1(20,11)            <= s_out1(21,11);
	s_in2(20,11)            <= s_out2(21,12);
	s_locks_lower_in(20,11) <= s_locks_lower_out(21,11);

		normal_cell_20_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,12),
			fetch              => s_fetch(20,12),
			data_in            => s_data_in(20,12),
			data_out           => s_data_out(20,12),
			out1               => s_out1(20,12),
			out2               => s_out2(20,12),
			lock_lower_row_out => s_locks_lower_out(20,12),
			lock_lower_row_in  => s_locks_lower_in(20,12),
			in1                => s_in1(20,12),
			in2                => s_in2(20,12),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(12)
		);
	s_in1(20,12)            <= s_out1(21,12);
	s_in2(20,12)            <= s_out2(21,13);
	s_locks_lower_in(20,12) <= s_locks_lower_out(21,12);

		normal_cell_20_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,13),
			fetch              => s_fetch(20,13),
			data_in            => s_data_in(20,13),
			data_out           => s_data_out(20,13),
			out1               => s_out1(20,13),
			out2               => s_out2(20,13),
			lock_lower_row_out => s_locks_lower_out(20,13),
			lock_lower_row_in  => s_locks_lower_in(20,13),
			in1                => s_in1(20,13),
			in2                => s_in2(20,13),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(13)
		);
	s_in1(20,13)            <= s_out1(21,13);
	s_in2(20,13)            <= s_out2(21,14);
	s_locks_lower_in(20,13) <= s_locks_lower_out(21,13);

		normal_cell_20_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,14),
			fetch              => s_fetch(20,14),
			data_in            => s_data_in(20,14),
			data_out           => s_data_out(20,14),
			out1               => s_out1(20,14),
			out2               => s_out2(20,14),
			lock_lower_row_out => s_locks_lower_out(20,14),
			lock_lower_row_in  => s_locks_lower_in(20,14),
			in1                => s_in1(20,14),
			in2                => s_in2(20,14),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(14)
		);
	s_in1(20,14)            <= s_out1(21,14);
	s_in2(20,14)            <= s_out2(21,15);
	s_locks_lower_in(20,14) <= s_locks_lower_out(21,14);

		normal_cell_20_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,15),
			fetch              => s_fetch(20,15),
			data_in            => s_data_in(20,15),
			data_out           => s_data_out(20,15),
			out1               => s_out1(20,15),
			out2               => s_out2(20,15),
			lock_lower_row_out => s_locks_lower_out(20,15),
			lock_lower_row_in  => s_locks_lower_in(20,15),
			in1                => s_in1(20,15),
			in2                => s_in2(20,15),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(15)
		);
	s_in1(20,15)            <= s_out1(21,15);
	s_in2(20,15)            <= s_out2(21,16);
	s_locks_lower_in(20,15) <= s_locks_lower_out(21,15);

		normal_cell_20_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,16),
			fetch              => s_fetch(20,16),
			data_in            => s_data_in(20,16),
			data_out           => s_data_out(20,16),
			out1               => s_out1(20,16),
			out2               => s_out2(20,16),
			lock_lower_row_out => s_locks_lower_out(20,16),
			lock_lower_row_in  => s_locks_lower_in(20,16),
			in1                => s_in1(20,16),
			in2                => s_in2(20,16),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(16)
		);
	s_in1(20,16)            <= s_out1(21,16);
	s_in2(20,16)            <= s_out2(21,17);
	s_locks_lower_in(20,16) <= s_locks_lower_out(21,16);

		normal_cell_20_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,17),
			fetch              => s_fetch(20,17),
			data_in            => s_data_in(20,17),
			data_out           => s_data_out(20,17),
			out1               => s_out1(20,17),
			out2               => s_out2(20,17),
			lock_lower_row_out => s_locks_lower_out(20,17),
			lock_lower_row_in  => s_locks_lower_in(20,17),
			in1                => s_in1(20,17),
			in2                => s_in2(20,17),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(17)
		);
	s_in1(20,17)            <= s_out1(21,17);
	s_in2(20,17)            <= s_out2(21,18);
	s_locks_lower_in(20,17) <= s_locks_lower_out(21,17);

		normal_cell_20_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,18),
			fetch              => s_fetch(20,18),
			data_in            => s_data_in(20,18),
			data_out           => s_data_out(20,18),
			out1               => s_out1(20,18),
			out2               => s_out2(20,18),
			lock_lower_row_out => s_locks_lower_out(20,18),
			lock_lower_row_in  => s_locks_lower_in(20,18),
			in1                => s_in1(20,18),
			in2                => s_in2(20,18),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(18)
		);
	s_in1(20,18)            <= s_out1(21,18);
	s_in2(20,18)            <= s_out2(21,19);
	s_locks_lower_in(20,18) <= s_locks_lower_out(21,18);

		normal_cell_20_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,19),
			fetch              => s_fetch(20,19),
			data_in            => s_data_in(20,19),
			data_out           => s_data_out(20,19),
			out1               => s_out1(20,19),
			out2               => s_out2(20,19),
			lock_lower_row_out => s_locks_lower_out(20,19),
			lock_lower_row_in  => s_locks_lower_in(20,19),
			in1                => s_in1(20,19),
			in2                => s_in2(20,19),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(19)
		);
	s_in1(20,19)            <= s_out1(21,19);
	s_in2(20,19)            <= s_out2(21,20);
	s_locks_lower_in(20,19) <= s_locks_lower_out(21,19);

		normal_cell_20_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,20),
			fetch              => s_fetch(20,20),
			data_in            => s_data_in(20,20),
			data_out           => s_data_out(20,20),
			out1               => s_out1(20,20),
			out2               => s_out2(20,20),
			lock_lower_row_out => s_locks_lower_out(20,20),
			lock_lower_row_in  => s_locks_lower_in(20,20),
			in1                => s_in1(20,20),
			in2                => s_in2(20,20),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(20)
		);
	s_in1(20,20)            <= s_out1(21,20);
	s_in2(20,20)            <= s_out2(21,21);
	s_locks_lower_in(20,20) <= s_locks_lower_out(21,20);

		normal_cell_20_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,21),
			fetch              => s_fetch(20,21),
			data_in            => s_data_in(20,21),
			data_out           => s_data_out(20,21),
			out1               => s_out1(20,21),
			out2               => s_out2(20,21),
			lock_lower_row_out => s_locks_lower_out(20,21),
			lock_lower_row_in  => s_locks_lower_in(20,21),
			in1                => s_in1(20,21),
			in2                => s_in2(20,21),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(21)
		);
	s_in1(20,21)            <= s_out1(21,21);
	s_in2(20,21)            <= s_out2(21,22);
	s_locks_lower_in(20,21) <= s_locks_lower_out(21,21);

		normal_cell_20_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,22),
			fetch              => s_fetch(20,22),
			data_in            => s_data_in(20,22),
			data_out           => s_data_out(20,22),
			out1               => s_out1(20,22),
			out2               => s_out2(20,22),
			lock_lower_row_out => s_locks_lower_out(20,22),
			lock_lower_row_in  => s_locks_lower_in(20,22),
			in1                => s_in1(20,22),
			in2                => s_in2(20,22),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(22)
		);
	s_in1(20,22)            <= s_out1(21,22);
	s_in2(20,22)            <= s_out2(21,23);
	s_locks_lower_in(20,22) <= s_locks_lower_out(21,22);

		normal_cell_20_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,23),
			fetch              => s_fetch(20,23),
			data_in            => s_data_in(20,23),
			data_out           => s_data_out(20,23),
			out1               => s_out1(20,23),
			out2               => s_out2(20,23),
			lock_lower_row_out => s_locks_lower_out(20,23),
			lock_lower_row_in  => s_locks_lower_in(20,23),
			in1                => s_in1(20,23),
			in2                => s_in2(20,23),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(23)
		);
	s_in1(20,23)            <= s_out1(21,23);
	s_in2(20,23)            <= s_out2(21,24);
	s_locks_lower_in(20,23) <= s_locks_lower_out(21,23);

		normal_cell_20_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,24),
			fetch              => s_fetch(20,24),
			data_in            => s_data_in(20,24),
			data_out           => s_data_out(20,24),
			out1               => s_out1(20,24),
			out2               => s_out2(20,24),
			lock_lower_row_out => s_locks_lower_out(20,24),
			lock_lower_row_in  => s_locks_lower_in(20,24),
			in1                => s_in1(20,24),
			in2                => s_in2(20,24),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(24)
		);
	s_in1(20,24)            <= s_out1(21,24);
	s_in2(20,24)            <= s_out2(21,25);
	s_locks_lower_in(20,24) <= s_locks_lower_out(21,24);

		normal_cell_20_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,25),
			fetch              => s_fetch(20,25),
			data_in            => s_data_in(20,25),
			data_out           => s_data_out(20,25),
			out1               => s_out1(20,25),
			out2               => s_out2(20,25),
			lock_lower_row_out => s_locks_lower_out(20,25),
			lock_lower_row_in  => s_locks_lower_in(20,25),
			in1                => s_in1(20,25),
			in2                => s_in2(20,25),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(25)
		);
	s_in1(20,25)            <= s_out1(21,25);
	s_in2(20,25)            <= s_out2(21,26);
	s_locks_lower_in(20,25) <= s_locks_lower_out(21,25);

		normal_cell_20_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,26),
			fetch              => s_fetch(20,26),
			data_in            => s_data_in(20,26),
			data_out           => s_data_out(20,26),
			out1               => s_out1(20,26),
			out2               => s_out2(20,26),
			lock_lower_row_out => s_locks_lower_out(20,26),
			lock_lower_row_in  => s_locks_lower_in(20,26),
			in1                => s_in1(20,26),
			in2                => s_in2(20,26),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(26)
		);
	s_in1(20,26)            <= s_out1(21,26);
	s_in2(20,26)            <= s_out2(21,27);
	s_locks_lower_in(20,26) <= s_locks_lower_out(21,26);

		normal_cell_20_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,27),
			fetch              => s_fetch(20,27),
			data_in            => s_data_in(20,27),
			data_out           => s_data_out(20,27),
			out1               => s_out1(20,27),
			out2               => s_out2(20,27),
			lock_lower_row_out => s_locks_lower_out(20,27),
			lock_lower_row_in  => s_locks_lower_in(20,27),
			in1                => s_in1(20,27),
			in2                => s_in2(20,27),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(27)
		);
	s_in1(20,27)            <= s_out1(21,27);
	s_in2(20,27)            <= s_out2(21,28);
	s_locks_lower_in(20,27) <= s_locks_lower_out(21,27);

		normal_cell_20_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,28),
			fetch              => s_fetch(20,28),
			data_in            => s_data_in(20,28),
			data_out           => s_data_out(20,28),
			out1               => s_out1(20,28),
			out2               => s_out2(20,28),
			lock_lower_row_out => s_locks_lower_out(20,28),
			lock_lower_row_in  => s_locks_lower_in(20,28),
			in1                => s_in1(20,28),
			in2                => s_in2(20,28),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(28)
		);
	s_in1(20,28)            <= s_out1(21,28);
	s_in2(20,28)            <= s_out2(21,29);
	s_locks_lower_in(20,28) <= s_locks_lower_out(21,28);

		normal_cell_20_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,29),
			fetch              => s_fetch(20,29),
			data_in            => s_data_in(20,29),
			data_out           => s_data_out(20,29),
			out1               => s_out1(20,29),
			out2               => s_out2(20,29),
			lock_lower_row_out => s_locks_lower_out(20,29),
			lock_lower_row_in  => s_locks_lower_in(20,29),
			in1                => s_in1(20,29),
			in2                => s_in2(20,29),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(29)
		);
	s_in1(20,29)            <= s_out1(21,29);
	s_in2(20,29)            <= s_out2(21,30);
	s_locks_lower_in(20,29) <= s_locks_lower_out(21,29);

		normal_cell_20_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,30),
			fetch              => s_fetch(20,30),
			data_in            => s_data_in(20,30),
			data_out           => s_data_out(20,30),
			out1               => s_out1(20,30),
			out2               => s_out2(20,30),
			lock_lower_row_out => s_locks_lower_out(20,30),
			lock_lower_row_in  => s_locks_lower_in(20,30),
			in1                => s_in1(20,30),
			in2                => s_in2(20,30),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(30)
		);
	s_in1(20,30)            <= s_out1(21,30);
	s_in2(20,30)            <= s_out2(21,31);
	s_locks_lower_in(20,30) <= s_locks_lower_out(21,30);

		normal_cell_20_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,31),
			fetch              => s_fetch(20,31),
			data_in            => s_data_in(20,31),
			data_out           => s_data_out(20,31),
			out1               => s_out1(20,31),
			out2               => s_out2(20,31),
			lock_lower_row_out => s_locks_lower_out(20,31),
			lock_lower_row_in  => s_locks_lower_in(20,31),
			in1                => s_in1(20,31),
			in2                => s_in2(20,31),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(31)
		);
	s_in1(20,31)            <= s_out1(21,31);
	s_in2(20,31)            <= s_out2(21,32);
	s_locks_lower_in(20,31) <= s_locks_lower_out(21,31);

		normal_cell_20_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,32),
			fetch              => s_fetch(20,32),
			data_in            => s_data_in(20,32),
			data_out           => s_data_out(20,32),
			out1               => s_out1(20,32),
			out2               => s_out2(20,32),
			lock_lower_row_out => s_locks_lower_out(20,32),
			lock_lower_row_in  => s_locks_lower_in(20,32),
			in1                => s_in1(20,32),
			in2                => s_in2(20,32),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(32)
		);
	s_in1(20,32)            <= s_out1(21,32);
	s_in2(20,32)            <= s_out2(21,33);
	s_locks_lower_in(20,32) <= s_locks_lower_out(21,32);

		normal_cell_20_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,33),
			fetch              => s_fetch(20,33),
			data_in            => s_data_in(20,33),
			data_out           => s_data_out(20,33),
			out1               => s_out1(20,33),
			out2               => s_out2(20,33),
			lock_lower_row_out => s_locks_lower_out(20,33),
			lock_lower_row_in  => s_locks_lower_in(20,33),
			in1                => s_in1(20,33),
			in2                => s_in2(20,33),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(33)
		);
	s_in1(20,33)            <= s_out1(21,33);
	s_in2(20,33)            <= s_out2(21,34);
	s_locks_lower_in(20,33) <= s_locks_lower_out(21,33);

		normal_cell_20_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,34),
			fetch              => s_fetch(20,34),
			data_in            => s_data_in(20,34),
			data_out           => s_data_out(20,34),
			out1               => s_out1(20,34),
			out2               => s_out2(20,34),
			lock_lower_row_out => s_locks_lower_out(20,34),
			lock_lower_row_in  => s_locks_lower_in(20,34),
			in1                => s_in1(20,34),
			in2                => s_in2(20,34),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(34)
		);
	s_in1(20,34)            <= s_out1(21,34);
	s_in2(20,34)            <= s_out2(21,35);
	s_locks_lower_in(20,34) <= s_locks_lower_out(21,34);

		normal_cell_20_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,35),
			fetch              => s_fetch(20,35),
			data_in            => s_data_in(20,35),
			data_out           => s_data_out(20,35),
			out1               => s_out1(20,35),
			out2               => s_out2(20,35),
			lock_lower_row_out => s_locks_lower_out(20,35),
			lock_lower_row_in  => s_locks_lower_in(20,35),
			in1                => s_in1(20,35),
			in2                => s_in2(20,35),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(35)
		);
	s_in1(20,35)            <= s_out1(21,35);
	s_in2(20,35)            <= s_out2(21,36);
	s_locks_lower_in(20,35) <= s_locks_lower_out(21,35);

		normal_cell_20_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,36),
			fetch              => s_fetch(20,36),
			data_in            => s_data_in(20,36),
			data_out           => s_data_out(20,36),
			out1               => s_out1(20,36),
			out2               => s_out2(20,36),
			lock_lower_row_out => s_locks_lower_out(20,36),
			lock_lower_row_in  => s_locks_lower_in(20,36),
			in1                => s_in1(20,36),
			in2                => s_in2(20,36),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(36)
		);
	s_in1(20,36)            <= s_out1(21,36);
	s_in2(20,36)            <= s_out2(21,37);
	s_locks_lower_in(20,36) <= s_locks_lower_out(21,36);

		normal_cell_20_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,37),
			fetch              => s_fetch(20,37),
			data_in            => s_data_in(20,37),
			data_out           => s_data_out(20,37),
			out1               => s_out1(20,37),
			out2               => s_out2(20,37),
			lock_lower_row_out => s_locks_lower_out(20,37),
			lock_lower_row_in  => s_locks_lower_in(20,37),
			in1                => s_in1(20,37),
			in2                => s_in2(20,37),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(37)
		);
	s_in1(20,37)            <= s_out1(21,37);
	s_in2(20,37)            <= s_out2(21,38);
	s_locks_lower_in(20,37) <= s_locks_lower_out(21,37);

		normal_cell_20_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,38),
			fetch              => s_fetch(20,38),
			data_in            => s_data_in(20,38),
			data_out           => s_data_out(20,38),
			out1               => s_out1(20,38),
			out2               => s_out2(20,38),
			lock_lower_row_out => s_locks_lower_out(20,38),
			lock_lower_row_in  => s_locks_lower_in(20,38),
			in1                => s_in1(20,38),
			in2                => s_in2(20,38),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(38)
		);
	s_in1(20,38)            <= s_out1(21,38);
	s_in2(20,38)            <= s_out2(21,39);
	s_locks_lower_in(20,38) <= s_locks_lower_out(21,38);

		normal_cell_20_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,39),
			fetch              => s_fetch(20,39),
			data_in            => s_data_in(20,39),
			data_out           => s_data_out(20,39),
			out1               => s_out1(20,39),
			out2               => s_out2(20,39),
			lock_lower_row_out => s_locks_lower_out(20,39),
			lock_lower_row_in  => s_locks_lower_in(20,39),
			in1                => s_in1(20,39),
			in2                => s_in2(20,39),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(39)
		);
	s_in1(20,39)            <= s_out1(21,39);
	s_in2(20,39)            <= s_out2(21,40);
	s_locks_lower_in(20,39) <= s_locks_lower_out(21,39);

		normal_cell_20_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,40),
			fetch              => s_fetch(20,40),
			data_in            => s_data_in(20,40),
			data_out           => s_data_out(20,40),
			out1               => s_out1(20,40),
			out2               => s_out2(20,40),
			lock_lower_row_out => s_locks_lower_out(20,40),
			lock_lower_row_in  => s_locks_lower_in(20,40),
			in1                => s_in1(20,40),
			in2                => s_in2(20,40),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(40)
		);
	s_in1(20,40)            <= s_out1(21,40);
	s_in2(20,40)            <= s_out2(21,41);
	s_locks_lower_in(20,40) <= s_locks_lower_out(21,40);

		normal_cell_20_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,41),
			fetch              => s_fetch(20,41),
			data_in            => s_data_in(20,41),
			data_out           => s_data_out(20,41),
			out1               => s_out1(20,41),
			out2               => s_out2(20,41),
			lock_lower_row_out => s_locks_lower_out(20,41),
			lock_lower_row_in  => s_locks_lower_in(20,41),
			in1                => s_in1(20,41),
			in2                => s_in2(20,41),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(41)
		);
	s_in1(20,41)            <= s_out1(21,41);
	s_in2(20,41)            <= s_out2(21,42);
	s_locks_lower_in(20,41) <= s_locks_lower_out(21,41);

		normal_cell_20_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,42),
			fetch              => s_fetch(20,42),
			data_in            => s_data_in(20,42),
			data_out           => s_data_out(20,42),
			out1               => s_out1(20,42),
			out2               => s_out2(20,42),
			lock_lower_row_out => s_locks_lower_out(20,42),
			lock_lower_row_in  => s_locks_lower_in(20,42),
			in1                => s_in1(20,42),
			in2                => s_in2(20,42),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(42)
		);
	s_in1(20,42)            <= s_out1(21,42);
	s_in2(20,42)            <= s_out2(21,43);
	s_locks_lower_in(20,42) <= s_locks_lower_out(21,42);

		normal_cell_20_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,43),
			fetch              => s_fetch(20,43),
			data_in            => s_data_in(20,43),
			data_out           => s_data_out(20,43),
			out1               => s_out1(20,43),
			out2               => s_out2(20,43),
			lock_lower_row_out => s_locks_lower_out(20,43),
			lock_lower_row_in  => s_locks_lower_in(20,43),
			in1                => s_in1(20,43),
			in2                => s_in2(20,43),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(43)
		);
	s_in1(20,43)            <= s_out1(21,43);
	s_in2(20,43)            <= s_out2(21,44);
	s_locks_lower_in(20,43) <= s_locks_lower_out(21,43);

		normal_cell_20_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,44),
			fetch              => s_fetch(20,44),
			data_in            => s_data_in(20,44),
			data_out           => s_data_out(20,44),
			out1               => s_out1(20,44),
			out2               => s_out2(20,44),
			lock_lower_row_out => s_locks_lower_out(20,44),
			lock_lower_row_in  => s_locks_lower_in(20,44),
			in1                => s_in1(20,44),
			in2                => s_in2(20,44),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(44)
		);
	s_in1(20,44)            <= s_out1(21,44);
	s_in2(20,44)            <= s_out2(21,45);
	s_locks_lower_in(20,44) <= s_locks_lower_out(21,44);

		normal_cell_20_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,45),
			fetch              => s_fetch(20,45),
			data_in            => s_data_in(20,45),
			data_out           => s_data_out(20,45),
			out1               => s_out1(20,45),
			out2               => s_out2(20,45),
			lock_lower_row_out => s_locks_lower_out(20,45),
			lock_lower_row_in  => s_locks_lower_in(20,45),
			in1                => s_in1(20,45),
			in2                => s_in2(20,45),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(45)
		);
	s_in1(20,45)            <= s_out1(21,45);
	s_in2(20,45)            <= s_out2(21,46);
	s_locks_lower_in(20,45) <= s_locks_lower_out(21,45);

		normal_cell_20_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,46),
			fetch              => s_fetch(20,46),
			data_in            => s_data_in(20,46),
			data_out           => s_data_out(20,46),
			out1               => s_out1(20,46),
			out2               => s_out2(20,46),
			lock_lower_row_out => s_locks_lower_out(20,46),
			lock_lower_row_in  => s_locks_lower_in(20,46),
			in1                => s_in1(20,46),
			in2                => s_in2(20,46),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(46)
		);
	s_in1(20,46)            <= s_out1(21,46);
	s_in2(20,46)            <= s_out2(21,47);
	s_locks_lower_in(20,46) <= s_locks_lower_out(21,46);

		normal_cell_20_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,47),
			fetch              => s_fetch(20,47),
			data_in            => s_data_in(20,47),
			data_out           => s_data_out(20,47),
			out1               => s_out1(20,47),
			out2               => s_out2(20,47),
			lock_lower_row_out => s_locks_lower_out(20,47),
			lock_lower_row_in  => s_locks_lower_in(20,47),
			in1                => s_in1(20,47),
			in2                => s_in2(20,47),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(47)
		);
	s_in1(20,47)            <= s_out1(21,47);
	s_in2(20,47)            <= s_out2(21,48);
	s_locks_lower_in(20,47) <= s_locks_lower_out(21,47);

		normal_cell_20_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,48),
			fetch              => s_fetch(20,48),
			data_in            => s_data_in(20,48),
			data_out           => s_data_out(20,48),
			out1               => s_out1(20,48),
			out2               => s_out2(20,48),
			lock_lower_row_out => s_locks_lower_out(20,48),
			lock_lower_row_in  => s_locks_lower_in(20,48),
			in1                => s_in1(20,48),
			in2                => s_in2(20,48),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(48)
		);
	s_in1(20,48)            <= s_out1(21,48);
	s_in2(20,48)            <= s_out2(21,49);
	s_locks_lower_in(20,48) <= s_locks_lower_out(21,48);

		normal_cell_20_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,49),
			fetch              => s_fetch(20,49),
			data_in            => s_data_in(20,49),
			data_out           => s_data_out(20,49),
			out1               => s_out1(20,49),
			out2               => s_out2(20,49),
			lock_lower_row_out => s_locks_lower_out(20,49),
			lock_lower_row_in  => s_locks_lower_in(20,49),
			in1                => s_in1(20,49),
			in2                => s_in2(20,49),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(49)
		);
	s_in1(20,49)            <= s_out1(21,49);
	s_in2(20,49)            <= s_out2(21,50);
	s_locks_lower_in(20,49) <= s_locks_lower_out(21,49);

		normal_cell_20_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,50),
			fetch              => s_fetch(20,50),
			data_in            => s_data_in(20,50),
			data_out           => s_data_out(20,50),
			out1               => s_out1(20,50),
			out2               => s_out2(20,50),
			lock_lower_row_out => s_locks_lower_out(20,50),
			lock_lower_row_in  => s_locks_lower_in(20,50),
			in1                => s_in1(20,50),
			in2                => s_in2(20,50),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(50)
		);
	s_in1(20,50)            <= s_out1(21,50);
	s_in2(20,50)            <= s_out2(21,51);
	s_locks_lower_in(20,50) <= s_locks_lower_out(21,50);

		normal_cell_20_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,51),
			fetch              => s_fetch(20,51),
			data_in            => s_data_in(20,51),
			data_out           => s_data_out(20,51),
			out1               => s_out1(20,51),
			out2               => s_out2(20,51),
			lock_lower_row_out => s_locks_lower_out(20,51),
			lock_lower_row_in  => s_locks_lower_in(20,51),
			in1                => s_in1(20,51),
			in2                => s_in2(20,51),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(51)
		);
	s_in1(20,51)            <= s_out1(21,51);
	s_in2(20,51)            <= s_out2(21,52);
	s_locks_lower_in(20,51) <= s_locks_lower_out(21,51);

		normal_cell_20_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,52),
			fetch              => s_fetch(20,52),
			data_in            => s_data_in(20,52),
			data_out           => s_data_out(20,52),
			out1               => s_out1(20,52),
			out2               => s_out2(20,52),
			lock_lower_row_out => s_locks_lower_out(20,52),
			lock_lower_row_in  => s_locks_lower_in(20,52),
			in1                => s_in1(20,52),
			in2                => s_in2(20,52),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(52)
		);
	s_in1(20,52)            <= s_out1(21,52);
	s_in2(20,52)            <= s_out2(21,53);
	s_locks_lower_in(20,52) <= s_locks_lower_out(21,52);

		normal_cell_20_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,53),
			fetch              => s_fetch(20,53),
			data_in            => s_data_in(20,53),
			data_out           => s_data_out(20,53),
			out1               => s_out1(20,53),
			out2               => s_out2(20,53),
			lock_lower_row_out => s_locks_lower_out(20,53),
			lock_lower_row_in  => s_locks_lower_in(20,53),
			in1                => s_in1(20,53),
			in2                => s_in2(20,53),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(53)
		);
	s_in1(20,53)            <= s_out1(21,53);
	s_in2(20,53)            <= s_out2(21,54);
	s_locks_lower_in(20,53) <= s_locks_lower_out(21,53);

		normal_cell_20_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,54),
			fetch              => s_fetch(20,54),
			data_in            => s_data_in(20,54),
			data_out           => s_data_out(20,54),
			out1               => s_out1(20,54),
			out2               => s_out2(20,54),
			lock_lower_row_out => s_locks_lower_out(20,54),
			lock_lower_row_in  => s_locks_lower_in(20,54),
			in1                => s_in1(20,54),
			in2                => s_in2(20,54),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(54)
		);
	s_in1(20,54)            <= s_out1(21,54);
	s_in2(20,54)            <= s_out2(21,55);
	s_locks_lower_in(20,54) <= s_locks_lower_out(21,54);

		normal_cell_20_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,55),
			fetch              => s_fetch(20,55),
			data_in            => s_data_in(20,55),
			data_out           => s_data_out(20,55),
			out1               => s_out1(20,55),
			out2               => s_out2(20,55),
			lock_lower_row_out => s_locks_lower_out(20,55),
			lock_lower_row_in  => s_locks_lower_in(20,55),
			in1                => s_in1(20,55),
			in2                => s_in2(20,55),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(55)
		);
	s_in1(20,55)            <= s_out1(21,55);
	s_in2(20,55)            <= s_out2(21,56);
	s_locks_lower_in(20,55) <= s_locks_lower_out(21,55);

		normal_cell_20_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,56),
			fetch              => s_fetch(20,56),
			data_in            => s_data_in(20,56),
			data_out           => s_data_out(20,56),
			out1               => s_out1(20,56),
			out2               => s_out2(20,56),
			lock_lower_row_out => s_locks_lower_out(20,56),
			lock_lower_row_in  => s_locks_lower_in(20,56),
			in1                => s_in1(20,56),
			in2                => s_in2(20,56),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(56)
		);
	s_in1(20,56)            <= s_out1(21,56);
	s_in2(20,56)            <= s_out2(21,57);
	s_locks_lower_in(20,56) <= s_locks_lower_out(21,56);

		normal_cell_20_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,57),
			fetch              => s_fetch(20,57),
			data_in            => s_data_in(20,57),
			data_out           => s_data_out(20,57),
			out1               => s_out1(20,57),
			out2               => s_out2(20,57),
			lock_lower_row_out => s_locks_lower_out(20,57),
			lock_lower_row_in  => s_locks_lower_in(20,57),
			in1                => s_in1(20,57),
			in2                => s_in2(20,57),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(57)
		);
	s_in1(20,57)            <= s_out1(21,57);
	s_in2(20,57)            <= s_out2(21,58);
	s_locks_lower_in(20,57) <= s_locks_lower_out(21,57);

		normal_cell_20_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,58),
			fetch              => s_fetch(20,58),
			data_in            => s_data_in(20,58),
			data_out           => s_data_out(20,58),
			out1               => s_out1(20,58),
			out2               => s_out2(20,58),
			lock_lower_row_out => s_locks_lower_out(20,58),
			lock_lower_row_in  => s_locks_lower_in(20,58),
			in1                => s_in1(20,58),
			in2                => s_in2(20,58),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(58)
		);
	s_in1(20,58)            <= s_out1(21,58);
	s_in2(20,58)            <= s_out2(21,59);
	s_locks_lower_in(20,58) <= s_locks_lower_out(21,58);

		normal_cell_20_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,59),
			fetch              => s_fetch(20,59),
			data_in            => s_data_in(20,59),
			data_out           => s_data_out(20,59),
			out1               => s_out1(20,59),
			out2               => s_out2(20,59),
			lock_lower_row_out => s_locks_lower_out(20,59),
			lock_lower_row_in  => s_locks_lower_in(20,59),
			in1                => s_in1(20,59),
			in2                => s_in2(20,59),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(59)
		);
	s_in1(20,59)            <= s_out1(21,59);
	s_in2(20,59)            <= s_out2(21,60);
	s_locks_lower_in(20,59) <= s_locks_lower_out(21,59);

		last_col_cell_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(20,60),
			fetch              => s_fetch(20,60),
			data_in            => s_data_in(20,60),
			data_out           => s_data_out(20,60),
			out1               => s_out1(20,60),
			out2               => s_out2(20,60),
			lock_lower_row_out => s_locks_lower_out(20,60),
			lock_lower_row_in  => s_locks_lower_in(20,60),
			in1                => s_in1(20,60),
			in2                => (others => '0'),
			lock_row           => s_locks(20),
			piv_found          => s_piv_found,
			row_data           => s_row_data(20),
			col_data           => s_col_data(60)
		);
	s_in1(20,60)            <= s_out1(21,60);
	s_locks_lower_in(20,60) <= s_locks_lower_out(21,60);

		normal_cell_21_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,1),
			fetch              => s_fetch(21,1),
			data_in            => s_data_in(21,1),
			data_out           => s_data_out(21,1),
			out1               => s_out1(21,1),
			out2               => s_out2(21,1),
			lock_lower_row_out => s_locks_lower_out(21,1),
			lock_lower_row_in  => s_locks_lower_in(21,1),
			in1                => s_in1(21,1),
			in2                => s_in2(21,1),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(1)
		);
	s_in1(21,1)            <= s_out1(22,1);
	s_in2(21,1)            <= s_out2(22,2);
	s_locks_lower_in(21,1) <= s_locks_lower_out(22,1);

		normal_cell_21_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,2),
			fetch              => s_fetch(21,2),
			data_in            => s_data_in(21,2),
			data_out           => s_data_out(21,2),
			out1               => s_out1(21,2),
			out2               => s_out2(21,2),
			lock_lower_row_out => s_locks_lower_out(21,2),
			lock_lower_row_in  => s_locks_lower_in(21,2),
			in1                => s_in1(21,2),
			in2                => s_in2(21,2),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(2)
		);
	s_in1(21,2)            <= s_out1(22,2);
	s_in2(21,2)            <= s_out2(22,3);
	s_locks_lower_in(21,2) <= s_locks_lower_out(22,2);

		normal_cell_21_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,3),
			fetch              => s_fetch(21,3),
			data_in            => s_data_in(21,3),
			data_out           => s_data_out(21,3),
			out1               => s_out1(21,3),
			out2               => s_out2(21,3),
			lock_lower_row_out => s_locks_lower_out(21,3),
			lock_lower_row_in  => s_locks_lower_in(21,3),
			in1                => s_in1(21,3),
			in2                => s_in2(21,3),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(3)
		);
	s_in1(21,3)            <= s_out1(22,3);
	s_in2(21,3)            <= s_out2(22,4);
	s_locks_lower_in(21,3) <= s_locks_lower_out(22,3);

		normal_cell_21_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,4),
			fetch              => s_fetch(21,4),
			data_in            => s_data_in(21,4),
			data_out           => s_data_out(21,4),
			out1               => s_out1(21,4),
			out2               => s_out2(21,4),
			lock_lower_row_out => s_locks_lower_out(21,4),
			lock_lower_row_in  => s_locks_lower_in(21,4),
			in1                => s_in1(21,4),
			in2                => s_in2(21,4),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(4)
		);
	s_in1(21,4)            <= s_out1(22,4);
	s_in2(21,4)            <= s_out2(22,5);
	s_locks_lower_in(21,4) <= s_locks_lower_out(22,4);

		normal_cell_21_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,5),
			fetch              => s_fetch(21,5),
			data_in            => s_data_in(21,5),
			data_out           => s_data_out(21,5),
			out1               => s_out1(21,5),
			out2               => s_out2(21,5),
			lock_lower_row_out => s_locks_lower_out(21,5),
			lock_lower_row_in  => s_locks_lower_in(21,5),
			in1                => s_in1(21,5),
			in2                => s_in2(21,5),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(5)
		);
	s_in1(21,5)            <= s_out1(22,5);
	s_in2(21,5)            <= s_out2(22,6);
	s_locks_lower_in(21,5) <= s_locks_lower_out(22,5);

		normal_cell_21_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,6),
			fetch              => s_fetch(21,6),
			data_in            => s_data_in(21,6),
			data_out           => s_data_out(21,6),
			out1               => s_out1(21,6),
			out2               => s_out2(21,6),
			lock_lower_row_out => s_locks_lower_out(21,6),
			lock_lower_row_in  => s_locks_lower_in(21,6),
			in1                => s_in1(21,6),
			in2                => s_in2(21,6),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(6)
		);
	s_in1(21,6)            <= s_out1(22,6);
	s_in2(21,6)            <= s_out2(22,7);
	s_locks_lower_in(21,6) <= s_locks_lower_out(22,6);

		normal_cell_21_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,7),
			fetch              => s_fetch(21,7),
			data_in            => s_data_in(21,7),
			data_out           => s_data_out(21,7),
			out1               => s_out1(21,7),
			out2               => s_out2(21,7),
			lock_lower_row_out => s_locks_lower_out(21,7),
			lock_lower_row_in  => s_locks_lower_in(21,7),
			in1                => s_in1(21,7),
			in2                => s_in2(21,7),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(7)
		);
	s_in1(21,7)            <= s_out1(22,7);
	s_in2(21,7)            <= s_out2(22,8);
	s_locks_lower_in(21,7) <= s_locks_lower_out(22,7);

		normal_cell_21_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,8),
			fetch              => s_fetch(21,8),
			data_in            => s_data_in(21,8),
			data_out           => s_data_out(21,8),
			out1               => s_out1(21,8),
			out2               => s_out2(21,8),
			lock_lower_row_out => s_locks_lower_out(21,8),
			lock_lower_row_in  => s_locks_lower_in(21,8),
			in1                => s_in1(21,8),
			in2                => s_in2(21,8),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(8)
		);
	s_in1(21,8)            <= s_out1(22,8);
	s_in2(21,8)            <= s_out2(22,9);
	s_locks_lower_in(21,8) <= s_locks_lower_out(22,8);

		normal_cell_21_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,9),
			fetch              => s_fetch(21,9),
			data_in            => s_data_in(21,9),
			data_out           => s_data_out(21,9),
			out1               => s_out1(21,9),
			out2               => s_out2(21,9),
			lock_lower_row_out => s_locks_lower_out(21,9),
			lock_lower_row_in  => s_locks_lower_in(21,9),
			in1                => s_in1(21,9),
			in2                => s_in2(21,9),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(9)
		);
	s_in1(21,9)            <= s_out1(22,9);
	s_in2(21,9)            <= s_out2(22,10);
	s_locks_lower_in(21,9) <= s_locks_lower_out(22,9);

		normal_cell_21_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,10),
			fetch              => s_fetch(21,10),
			data_in            => s_data_in(21,10),
			data_out           => s_data_out(21,10),
			out1               => s_out1(21,10),
			out2               => s_out2(21,10),
			lock_lower_row_out => s_locks_lower_out(21,10),
			lock_lower_row_in  => s_locks_lower_in(21,10),
			in1                => s_in1(21,10),
			in2                => s_in2(21,10),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(10)
		);
	s_in1(21,10)            <= s_out1(22,10);
	s_in2(21,10)            <= s_out2(22,11);
	s_locks_lower_in(21,10) <= s_locks_lower_out(22,10);

		normal_cell_21_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,11),
			fetch              => s_fetch(21,11),
			data_in            => s_data_in(21,11),
			data_out           => s_data_out(21,11),
			out1               => s_out1(21,11),
			out2               => s_out2(21,11),
			lock_lower_row_out => s_locks_lower_out(21,11),
			lock_lower_row_in  => s_locks_lower_in(21,11),
			in1                => s_in1(21,11),
			in2                => s_in2(21,11),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(11)
		);
	s_in1(21,11)            <= s_out1(22,11);
	s_in2(21,11)            <= s_out2(22,12);
	s_locks_lower_in(21,11) <= s_locks_lower_out(22,11);

		normal_cell_21_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,12),
			fetch              => s_fetch(21,12),
			data_in            => s_data_in(21,12),
			data_out           => s_data_out(21,12),
			out1               => s_out1(21,12),
			out2               => s_out2(21,12),
			lock_lower_row_out => s_locks_lower_out(21,12),
			lock_lower_row_in  => s_locks_lower_in(21,12),
			in1                => s_in1(21,12),
			in2                => s_in2(21,12),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(12)
		);
	s_in1(21,12)            <= s_out1(22,12);
	s_in2(21,12)            <= s_out2(22,13);
	s_locks_lower_in(21,12) <= s_locks_lower_out(22,12);

		normal_cell_21_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,13),
			fetch              => s_fetch(21,13),
			data_in            => s_data_in(21,13),
			data_out           => s_data_out(21,13),
			out1               => s_out1(21,13),
			out2               => s_out2(21,13),
			lock_lower_row_out => s_locks_lower_out(21,13),
			lock_lower_row_in  => s_locks_lower_in(21,13),
			in1                => s_in1(21,13),
			in2                => s_in2(21,13),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(13)
		);
	s_in1(21,13)            <= s_out1(22,13);
	s_in2(21,13)            <= s_out2(22,14);
	s_locks_lower_in(21,13) <= s_locks_lower_out(22,13);

		normal_cell_21_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,14),
			fetch              => s_fetch(21,14),
			data_in            => s_data_in(21,14),
			data_out           => s_data_out(21,14),
			out1               => s_out1(21,14),
			out2               => s_out2(21,14),
			lock_lower_row_out => s_locks_lower_out(21,14),
			lock_lower_row_in  => s_locks_lower_in(21,14),
			in1                => s_in1(21,14),
			in2                => s_in2(21,14),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(14)
		);
	s_in1(21,14)            <= s_out1(22,14);
	s_in2(21,14)            <= s_out2(22,15);
	s_locks_lower_in(21,14) <= s_locks_lower_out(22,14);

		normal_cell_21_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,15),
			fetch              => s_fetch(21,15),
			data_in            => s_data_in(21,15),
			data_out           => s_data_out(21,15),
			out1               => s_out1(21,15),
			out2               => s_out2(21,15),
			lock_lower_row_out => s_locks_lower_out(21,15),
			lock_lower_row_in  => s_locks_lower_in(21,15),
			in1                => s_in1(21,15),
			in2                => s_in2(21,15),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(15)
		);
	s_in1(21,15)            <= s_out1(22,15);
	s_in2(21,15)            <= s_out2(22,16);
	s_locks_lower_in(21,15) <= s_locks_lower_out(22,15);

		normal_cell_21_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,16),
			fetch              => s_fetch(21,16),
			data_in            => s_data_in(21,16),
			data_out           => s_data_out(21,16),
			out1               => s_out1(21,16),
			out2               => s_out2(21,16),
			lock_lower_row_out => s_locks_lower_out(21,16),
			lock_lower_row_in  => s_locks_lower_in(21,16),
			in1                => s_in1(21,16),
			in2                => s_in2(21,16),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(16)
		);
	s_in1(21,16)            <= s_out1(22,16);
	s_in2(21,16)            <= s_out2(22,17);
	s_locks_lower_in(21,16) <= s_locks_lower_out(22,16);

		normal_cell_21_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,17),
			fetch              => s_fetch(21,17),
			data_in            => s_data_in(21,17),
			data_out           => s_data_out(21,17),
			out1               => s_out1(21,17),
			out2               => s_out2(21,17),
			lock_lower_row_out => s_locks_lower_out(21,17),
			lock_lower_row_in  => s_locks_lower_in(21,17),
			in1                => s_in1(21,17),
			in2                => s_in2(21,17),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(17)
		);
	s_in1(21,17)            <= s_out1(22,17);
	s_in2(21,17)            <= s_out2(22,18);
	s_locks_lower_in(21,17) <= s_locks_lower_out(22,17);

		normal_cell_21_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,18),
			fetch              => s_fetch(21,18),
			data_in            => s_data_in(21,18),
			data_out           => s_data_out(21,18),
			out1               => s_out1(21,18),
			out2               => s_out2(21,18),
			lock_lower_row_out => s_locks_lower_out(21,18),
			lock_lower_row_in  => s_locks_lower_in(21,18),
			in1                => s_in1(21,18),
			in2                => s_in2(21,18),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(18)
		);
	s_in1(21,18)            <= s_out1(22,18);
	s_in2(21,18)            <= s_out2(22,19);
	s_locks_lower_in(21,18) <= s_locks_lower_out(22,18);

		normal_cell_21_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,19),
			fetch              => s_fetch(21,19),
			data_in            => s_data_in(21,19),
			data_out           => s_data_out(21,19),
			out1               => s_out1(21,19),
			out2               => s_out2(21,19),
			lock_lower_row_out => s_locks_lower_out(21,19),
			lock_lower_row_in  => s_locks_lower_in(21,19),
			in1                => s_in1(21,19),
			in2                => s_in2(21,19),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(19)
		);
	s_in1(21,19)            <= s_out1(22,19);
	s_in2(21,19)            <= s_out2(22,20);
	s_locks_lower_in(21,19) <= s_locks_lower_out(22,19);

		normal_cell_21_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,20),
			fetch              => s_fetch(21,20),
			data_in            => s_data_in(21,20),
			data_out           => s_data_out(21,20),
			out1               => s_out1(21,20),
			out2               => s_out2(21,20),
			lock_lower_row_out => s_locks_lower_out(21,20),
			lock_lower_row_in  => s_locks_lower_in(21,20),
			in1                => s_in1(21,20),
			in2                => s_in2(21,20),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(20)
		);
	s_in1(21,20)            <= s_out1(22,20);
	s_in2(21,20)            <= s_out2(22,21);
	s_locks_lower_in(21,20) <= s_locks_lower_out(22,20);

		normal_cell_21_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,21),
			fetch              => s_fetch(21,21),
			data_in            => s_data_in(21,21),
			data_out           => s_data_out(21,21),
			out1               => s_out1(21,21),
			out2               => s_out2(21,21),
			lock_lower_row_out => s_locks_lower_out(21,21),
			lock_lower_row_in  => s_locks_lower_in(21,21),
			in1                => s_in1(21,21),
			in2                => s_in2(21,21),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(21)
		);
	s_in1(21,21)            <= s_out1(22,21);
	s_in2(21,21)            <= s_out2(22,22);
	s_locks_lower_in(21,21) <= s_locks_lower_out(22,21);

		normal_cell_21_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,22),
			fetch              => s_fetch(21,22),
			data_in            => s_data_in(21,22),
			data_out           => s_data_out(21,22),
			out1               => s_out1(21,22),
			out2               => s_out2(21,22),
			lock_lower_row_out => s_locks_lower_out(21,22),
			lock_lower_row_in  => s_locks_lower_in(21,22),
			in1                => s_in1(21,22),
			in2                => s_in2(21,22),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(22)
		);
	s_in1(21,22)            <= s_out1(22,22);
	s_in2(21,22)            <= s_out2(22,23);
	s_locks_lower_in(21,22) <= s_locks_lower_out(22,22);

		normal_cell_21_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,23),
			fetch              => s_fetch(21,23),
			data_in            => s_data_in(21,23),
			data_out           => s_data_out(21,23),
			out1               => s_out1(21,23),
			out2               => s_out2(21,23),
			lock_lower_row_out => s_locks_lower_out(21,23),
			lock_lower_row_in  => s_locks_lower_in(21,23),
			in1                => s_in1(21,23),
			in2                => s_in2(21,23),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(23)
		);
	s_in1(21,23)            <= s_out1(22,23);
	s_in2(21,23)            <= s_out2(22,24);
	s_locks_lower_in(21,23) <= s_locks_lower_out(22,23);

		normal_cell_21_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,24),
			fetch              => s_fetch(21,24),
			data_in            => s_data_in(21,24),
			data_out           => s_data_out(21,24),
			out1               => s_out1(21,24),
			out2               => s_out2(21,24),
			lock_lower_row_out => s_locks_lower_out(21,24),
			lock_lower_row_in  => s_locks_lower_in(21,24),
			in1                => s_in1(21,24),
			in2                => s_in2(21,24),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(24)
		);
	s_in1(21,24)            <= s_out1(22,24);
	s_in2(21,24)            <= s_out2(22,25);
	s_locks_lower_in(21,24) <= s_locks_lower_out(22,24);

		normal_cell_21_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,25),
			fetch              => s_fetch(21,25),
			data_in            => s_data_in(21,25),
			data_out           => s_data_out(21,25),
			out1               => s_out1(21,25),
			out2               => s_out2(21,25),
			lock_lower_row_out => s_locks_lower_out(21,25),
			lock_lower_row_in  => s_locks_lower_in(21,25),
			in1                => s_in1(21,25),
			in2                => s_in2(21,25),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(25)
		);
	s_in1(21,25)            <= s_out1(22,25);
	s_in2(21,25)            <= s_out2(22,26);
	s_locks_lower_in(21,25) <= s_locks_lower_out(22,25);

		normal_cell_21_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,26),
			fetch              => s_fetch(21,26),
			data_in            => s_data_in(21,26),
			data_out           => s_data_out(21,26),
			out1               => s_out1(21,26),
			out2               => s_out2(21,26),
			lock_lower_row_out => s_locks_lower_out(21,26),
			lock_lower_row_in  => s_locks_lower_in(21,26),
			in1                => s_in1(21,26),
			in2                => s_in2(21,26),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(26)
		);
	s_in1(21,26)            <= s_out1(22,26);
	s_in2(21,26)            <= s_out2(22,27);
	s_locks_lower_in(21,26) <= s_locks_lower_out(22,26);

		normal_cell_21_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,27),
			fetch              => s_fetch(21,27),
			data_in            => s_data_in(21,27),
			data_out           => s_data_out(21,27),
			out1               => s_out1(21,27),
			out2               => s_out2(21,27),
			lock_lower_row_out => s_locks_lower_out(21,27),
			lock_lower_row_in  => s_locks_lower_in(21,27),
			in1                => s_in1(21,27),
			in2                => s_in2(21,27),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(27)
		);
	s_in1(21,27)            <= s_out1(22,27);
	s_in2(21,27)            <= s_out2(22,28);
	s_locks_lower_in(21,27) <= s_locks_lower_out(22,27);

		normal_cell_21_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,28),
			fetch              => s_fetch(21,28),
			data_in            => s_data_in(21,28),
			data_out           => s_data_out(21,28),
			out1               => s_out1(21,28),
			out2               => s_out2(21,28),
			lock_lower_row_out => s_locks_lower_out(21,28),
			lock_lower_row_in  => s_locks_lower_in(21,28),
			in1                => s_in1(21,28),
			in2                => s_in2(21,28),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(28)
		);
	s_in1(21,28)            <= s_out1(22,28);
	s_in2(21,28)            <= s_out2(22,29);
	s_locks_lower_in(21,28) <= s_locks_lower_out(22,28);

		normal_cell_21_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,29),
			fetch              => s_fetch(21,29),
			data_in            => s_data_in(21,29),
			data_out           => s_data_out(21,29),
			out1               => s_out1(21,29),
			out2               => s_out2(21,29),
			lock_lower_row_out => s_locks_lower_out(21,29),
			lock_lower_row_in  => s_locks_lower_in(21,29),
			in1                => s_in1(21,29),
			in2                => s_in2(21,29),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(29)
		);
	s_in1(21,29)            <= s_out1(22,29);
	s_in2(21,29)            <= s_out2(22,30);
	s_locks_lower_in(21,29) <= s_locks_lower_out(22,29);

		normal_cell_21_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,30),
			fetch              => s_fetch(21,30),
			data_in            => s_data_in(21,30),
			data_out           => s_data_out(21,30),
			out1               => s_out1(21,30),
			out2               => s_out2(21,30),
			lock_lower_row_out => s_locks_lower_out(21,30),
			lock_lower_row_in  => s_locks_lower_in(21,30),
			in1                => s_in1(21,30),
			in2                => s_in2(21,30),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(30)
		);
	s_in1(21,30)            <= s_out1(22,30);
	s_in2(21,30)            <= s_out2(22,31);
	s_locks_lower_in(21,30) <= s_locks_lower_out(22,30);

		normal_cell_21_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,31),
			fetch              => s_fetch(21,31),
			data_in            => s_data_in(21,31),
			data_out           => s_data_out(21,31),
			out1               => s_out1(21,31),
			out2               => s_out2(21,31),
			lock_lower_row_out => s_locks_lower_out(21,31),
			lock_lower_row_in  => s_locks_lower_in(21,31),
			in1                => s_in1(21,31),
			in2                => s_in2(21,31),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(31)
		);
	s_in1(21,31)            <= s_out1(22,31);
	s_in2(21,31)            <= s_out2(22,32);
	s_locks_lower_in(21,31) <= s_locks_lower_out(22,31);

		normal_cell_21_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,32),
			fetch              => s_fetch(21,32),
			data_in            => s_data_in(21,32),
			data_out           => s_data_out(21,32),
			out1               => s_out1(21,32),
			out2               => s_out2(21,32),
			lock_lower_row_out => s_locks_lower_out(21,32),
			lock_lower_row_in  => s_locks_lower_in(21,32),
			in1                => s_in1(21,32),
			in2                => s_in2(21,32),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(32)
		);
	s_in1(21,32)            <= s_out1(22,32);
	s_in2(21,32)            <= s_out2(22,33);
	s_locks_lower_in(21,32) <= s_locks_lower_out(22,32);

		normal_cell_21_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,33),
			fetch              => s_fetch(21,33),
			data_in            => s_data_in(21,33),
			data_out           => s_data_out(21,33),
			out1               => s_out1(21,33),
			out2               => s_out2(21,33),
			lock_lower_row_out => s_locks_lower_out(21,33),
			lock_lower_row_in  => s_locks_lower_in(21,33),
			in1                => s_in1(21,33),
			in2                => s_in2(21,33),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(33)
		);
	s_in1(21,33)            <= s_out1(22,33);
	s_in2(21,33)            <= s_out2(22,34);
	s_locks_lower_in(21,33) <= s_locks_lower_out(22,33);

		normal_cell_21_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,34),
			fetch              => s_fetch(21,34),
			data_in            => s_data_in(21,34),
			data_out           => s_data_out(21,34),
			out1               => s_out1(21,34),
			out2               => s_out2(21,34),
			lock_lower_row_out => s_locks_lower_out(21,34),
			lock_lower_row_in  => s_locks_lower_in(21,34),
			in1                => s_in1(21,34),
			in2                => s_in2(21,34),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(34)
		);
	s_in1(21,34)            <= s_out1(22,34);
	s_in2(21,34)            <= s_out2(22,35);
	s_locks_lower_in(21,34) <= s_locks_lower_out(22,34);

		normal_cell_21_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,35),
			fetch              => s_fetch(21,35),
			data_in            => s_data_in(21,35),
			data_out           => s_data_out(21,35),
			out1               => s_out1(21,35),
			out2               => s_out2(21,35),
			lock_lower_row_out => s_locks_lower_out(21,35),
			lock_lower_row_in  => s_locks_lower_in(21,35),
			in1                => s_in1(21,35),
			in2                => s_in2(21,35),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(35)
		);
	s_in1(21,35)            <= s_out1(22,35);
	s_in2(21,35)            <= s_out2(22,36);
	s_locks_lower_in(21,35) <= s_locks_lower_out(22,35);

		normal_cell_21_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,36),
			fetch              => s_fetch(21,36),
			data_in            => s_data_in(21,36),
			data_out           => s_data_out(21,36),
			out1               => s_out1(21,36),
			out2               => s_out2(21,36),
			lock_lower_row_out => s_locks_lower_out(21,36),
			lock_lower_row_in  => s_locks_lower_in(21,36),
			in1                => s_in1(21,36),
			in2                => s_in2(21,36),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(36)
		);
	s_in1(21,36)            <= s_out1(22,36);
	s_in2(21,36)            <= s_out2(22,37);
	s_locks_lower_in(21,36) <= s_locks_lower_out(22,36);

		normal_cell_21_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,37),
			fetch              => s_fetch(21,37),
			data_in            => s_data_in(21,37),
			data_out           => s_data_out(21,37),
			out1               => s_out1(21,37),
			out2               => s_out2(21,37),
			lock_lower_row_out => s_locks_lower_out(21,37),
			lock_lower_row_in  => s_locks_lower_in(21,37),
			in1                => s_in1(21,37),
			in2                => s_in2(21,37),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(37)
		);
	s_in1(21,37)            <= s_out1(22,37);
	s_in2(21,37)            <= s_out2(22,38);
	s_locks_lower_in(21,37) <= s_locks_lower_out(22,37);

		normal_cell_21_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,38),
			fetch              => s_fetch(21,38),
			data_in            => s_data_in(21,38),
			data_out           => s_data_out(21,38),
			out1               => s_out1(21,38),
			out2               => s_out2(21,38),
			lock_lower_row_out => s_locks_lower_out(21,38),
			lock_lower_row_in  => s_locks_lower_in(21,38),
			in1                => s_in1(21,38),
			in2                => s_in2(21,38),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(38)
		);
	s_in1(21,38)            <= s_out1(22,38);
	s_in2(21,38)            <= s_out2(22,39);
	s_locks_lower_in(21,38) <= s_locks_lower_out(22,38);

		normal_cell_21_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,39),
			fetch              => s_fetch(21,39),
			data_in            => s_data_in(21,39),
			data_out           => s_data_out(21,39),
			out1               => s_out1(21,39),
			out2               => s_out2(21,39),
			lock_lower_row_out => s_locks_lower_out(21,39),
			lock_lower_row_in  => s_locks_lower_in(21,39),
			in1                => s_in1(21,39),
			in2                => s_in2(21,39),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(39)
		);
	s_in1(21,39)            <= s_out1(22,39);
	s_in2(21,39)            <= s_out2(22,40);
	s_locks_lower_in(21,39) <= s_locks_lower_out(22,39);

		normal_cell_21_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,40),
			fetch              => s_fetch(21,40),
			data_in            => s_data_in(21,40),
			data_out           => s_data_out(21,40),
			out1               => s_out1(21,40),
			out2               => s_out2(21,40),
			lock_lower_row_out => s_locks_lower_out(21,40),
			lock_lower_row_in  => s_locks_lower_in(21,40),
			in1                => s_in1(21,40),
			in2                => s_in2(21,40),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(40)
		);
	s_in1(21,40)            <= s_out1(22,40);
	s_in2(21,40)            <= s_out2(22,41);
	s_locks_lower_in(21,40) <= s_locks_lower_out(22,40);

		normal_cell_21_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,41),
			fetch              => s_fetch(21,41),
			data_in            => s_data_in(21,41),
			data_out           => s_data_out(21,41),
			out1               => s_out1(21,41),
			out2               => s_out2(21,41),
			lock_lower_row_out => s_locks_lower_out(21,41),
			lock_lower_row_in  => s_locks_lower_in(21,41),
			in1                => s_in1(21,41),
			in2                => s_in2(21,41),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(41)
		);
	s_in1(21,41)            <= s_out1(22,41);
	s_in2(21,41)            <= s_out2(22,42);
	s_locks_lower_in(21,41) <= s_locks_lower_out(22,41);

		normal_cell_21_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,42),
			fetch              => s_fetch(21,42),
			data_in            => s_data_in(21,42),
			data_out           => s_data_out(21,42),
			out1               => s_out1(21,42),
			out2               => s_out2(21,42),
			lock_lower_row_out => s_locks_lower_out(21,42),
			lock_lower_row_in  => s_locks_lower_in(21,42),
			in1                => s_in1(21,42),
			in2                => s_in2(21,42),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(42)
		);
	s_in1(21,42)            <= s_out1(22,42);
	s_in2(21,42)            <= s_out2(22,43);
	s_locks_lower_in(21,42) <= s_locks_lower_out(22,42);

		normal_cell_21_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,43),
			fetch              => s_fetch(21,43),
			data_in            => s_data_in(21,43),
			data_out           => s_data_out(21,43),
			out1               => s_out1(21,43),
			out2               => s_out2(21,43),
			lock_lower_row_out => s_locks_lower_out(21,43),
			lock_lower_row_in  => s_locks_lower_in(21,43),
			in1                => s_in1(21,43),
			in2                => s_in2(21,43),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(43)
		);
	s_in1(21,43)            <= s_out1(22,43);
	s_in2(21,43)            <= s_out2(22,44);
	s_locks_lower_in(21,43) <= s_locks_lower_out(22,43);

		normal_cell_21_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,44),
			fetch              => s_fetch(21,44),
			data_in            => s_data_in(21,44),
			data_out           => s_data_out(21,44),
			out1               => s_out1(21,44),
			out2               => s_out2(21,44),
			lock_lower_row_out => s_locks_lower_out(21,44),
			lock_lower_row_in  => s_locks_lower_in(21,44),
			in1                => s_in1(21,44),
			in2                => s_in2(21,44),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(44)
		);
	s_in1(21,44)            <= s_out1(22,44);
	s_in2(21,44)            <= s_out2(22,45);
	s_locks_lower_in(21,44) <= s_locks_lower_out(22,44);

		normal_cell_21_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,45),
			fetch              => s_fetch(21,45),
			data_in            => s_data_in(21,45),
			data_out           => s_data_out(21,45),
			out1               => s_out1(21,45),
			out2               => s_out2(21,45),
			lock_lower_row_out => s_locks_lower_out(21,45),
			lock_lower_row_in  => s_locks_lower_in(21,45),
			in1                => s_in1(21,45),
			in2                => s_in2(21,45),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(45)
		);
	s_in1(21,45)            <= s_out1(22,45);
	s_in2(21,45)            <= s_out2(22,46);
	s_locks_lower_in(21,45) <= s_locks_lower_out(22,45);

		normal_cell_21_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,46),
			fetch              => s_fetch(21,46),
			data_in            => s_data_in(21,46),
			data_out           => s_data_out(21,46),
			out1               => s_out1(21,46),
			out2               => s_out2(21,46),
			lock_lower_row_out => s_locks_lower_out(21,46),
			lock_lower_row_in  => s_locks_lower_in(21,46),
			in1                => s_in1(21,46),
			in2                => s_in2(21,46),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(46)
		);
	s_in1(21,46)            <= s_out1(22,46);
	s_in2(21,46)            <= s_out2(22,47);
	s_locks_lower_in(21,46) <= s_locks_lower_out(22,46);

		normal_cell_21_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,47),
			fetch              => s_fetch(21,47),
			data_in            => s_data_in(21,47),
			data_out           => s_data_out(21,47),
			out1               => s_out1(21,47),
			out2               => s_out2(21,47),
			lock_lower_row_out => s_locks_lower_out(21,47),
			lock_lower_row_in  => s_locks_lower_in(21,47),
			in1                => s_in1(21,47),
			in2                => s_in2(21,47),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(47)
		);
	s_in1(21,47)            <= s_out1(22,47);
	s_in2(21,47)            <= s_out2(22,48);
	s_locks_lower_in(21,47) <= s_locks_lower_out(22,47);

		normal_cell_21_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,48),
			fetch              => s_fetch(21,48),
			data_in            => s_data_in(21,48),
			data_out           => s_data_out(21,48),
			out1               => s_out1(21,48),
			out2               => s_out2(21,48),
			lock_lower_row_out => s_locks_lower_out(21,48),
			lock_lower_row_in  => s_locks_lower_in(21,48),
			in1                => s_in1(21,48),
			in2                => s_in2(21,48),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(48)
		);
	s_in1(21,48)            <= s_out1(22,48);
	s_in2(21,48)            <= s_out2(22,49);
	s_locks_lower_in(21,48) <= s_locks_lower_out(22,48);

		normal_cell_21_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,49),
			fetch              => s_fetch(21,49),
			data_in            => s_data_in(21,49),
			data_out           => s_data_out(21,49),
			out1               => s_out1(21,49),
			out2               => s_out2(21,49),
			lock_lower_row_out => s_locks_lower_out(21,49),
			lock_lower_row_in  => s_locks_lower_in(21,49),
			in1                => s_in1(21,49),
			in2                => s_in2(21,49),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(49)
		);
	s_in1(21,49)            <= s_out1(22,49);
	s_in2(21,49)            <= s_out2(22,50);
	s_locks_lower_in(21,49) <= s_locks_lower_out(22,49);

		normal_cell_21_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,50),
			fetch              => s_fetch(21,50),
			data_in            => s_data_in(21,50),
			data_out           => s_data_out(21,50),
			out1               => s_out1(21,50),
			out2               => s_out2(21,50),
			lock_lower_row_out => s_locks_lower_out(21,50),
			lock_lower_row_in  => s_locks_lower_in(21,50),
			in1                => s_in1(21,50),
			in2                => s_in2(21,50),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(50)
		);
	s_in1(21,50)            <= s_out1(22,50);
	s_in2(21,50)            <= s_out2(22,51);
	s_locks_lower_in(21,50) <= s_locks_lower_out(22,50);

		normal_cell_21_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,51),
			fetch              => s_fetch(21,51),
			data_in            => s_data_in(21,51),
			data_out           => s_data_out(21,51),
			out1               => s_out1(21,51),
			out2               => s_out2(21,51),
			lock_lower_row_out => s_locks_lower_out(21,51),
			lock_lower_row_in  => s_locks_lower_in(21,51),
			in1                => s_in1(21,51),
			in2                => s_in2(21,51),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(51)
		);
	s_in1(21,51)            <= s_out1(22,51);
	s_in2(21,51)            <= s_out2(22,52);
	s_locks_lower_in(21,51) <= s_locks_lower_out(22,51);

		normal_cell_21_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,52),
			fetch              => s_fetch(21,52),
			data_in            => s_data_in(21,52),
			data_out           => s_data_out(21,52),
			out1               => s_out1(21,52),
			out2               => s_out2(21,52),
			lock_lower_row_out => s_locks_lower_out(21,52),
			lock_lower_row_in  => s_locks_lower_in(21,52),
			in1                => s_in1(21,52),
			in2                => s_in2(21,52),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(52)
		);
	s_in1(21,52)            <= s_out1(22,52);
	s_in2(21,52)            <= s_out2(22,53);
	s_locks_lower_in(21,52) <= s_locks_lower_out(22,52);

		normal_cell_21_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,53),
			fetch              => s_fetch(21,53),
			data_in            => s_data_in(21,53),
			data_out           => s_data_out(21,53),
			out1               => s_out1(21,53),
			out2               => s_out2(21,53),
			lock_lower_row_out => s_locks_lower_out(21,53),
			lock_lower_row_in  => s_locks_lower_in(21,53),
			in1                => s_in1(21,53),
			in2                => s_in2(21,53),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(53)
		);
	s_in1(21,53)            <= s_out1(22,53);
	s_in2(21,53)            <= s_out2(22,54);
	s_locks_lower_in(21,53) <= s_locks_lower_out(22,53);

		normal_cell_21_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,54),
			fetch              => s_fetch(21,54),
			data_in            => s_data_in(21,54),
			data_out           => s_data_out(21,54),
			out1               => s_out1(21,54),
			out2               => s_out2(21,54),
			lock_lower_row_out => s_locks_lower_out(21,54),
			lock_lower_row_in  => s_locks_lower_in(21,54),
			in1                => s_in1(21,54),
			in2                => s_in2(21,54),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(54)
		);
	s_in1(21,54)            <= s_out1(22,54);
	s_in2(21,54)            <= s_out2(22,55);
	s_locks_lower_in(21,54) <= s_locks_lower_out(22,54);

		normal_cell_21_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,55),
			fetch              => s_fetch(21,55),
			data_in            => s_data_in(21,55),
			data_out           => s_data_out(21,55),
			out1               => s_out1(21,55),
			out2               => s_out2(21,55),
			lock_lower_row_out => s_locks_lower_out(21,55),
			lock_lower_row_in  => s_locks_lower_in(21,55),
			in1                => s_in1(21,55),
			in2                => s_in2(21,55),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(55)
		);
	s_in1(21,55)            <= s_out1(22,55);
	s_in2(21,55)            <= s_out2(22,56);
	s_locks_lower_in(21,55) <= s_locks_lower_out(22,55);

		normal_cell_21_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,56),
			fetch              => s_fetch(21,56),
			data_in            => s_data_in(21,56),
			data_out           => s_data_out(21,56),
			out1               => s_out1(21,56),
			out2               => s_out2(21,56),
			lock_lower_row_out => s_locks_lower_out(21,56),
			lock_lower_row_in  => s_locks_lower_in(21,56),
			in1                => s_in1(21,56),
			in2                => s_in2(21,56),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(56)
		);
	s_in1(21,56)            <= s_out1(22,56);
	s_in2(21,56)            <= s_out2(22,57);
	s_locks_lower_in(21,56) <= s_locks_lower_out(22,56);

		normal_cell_21_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,57),
			fetch              => s_fetch(21,57),
			data_in            => s_data_in(21,57),
			data_out           => s_data_out(21,57),
			out1               => s_out1(21,57),
			out2               => s_out2(21,57),
			lock_lower_row_out => s_locks_lower_out(21,57),
			lock_lower_row_in  => s_locks_lower_in(21,57),
			in1                => s_in1(21,57),
			in2                => s_in2(21,57),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(57)
		);
	s_in1(21,57)            <= s_out1(22,57);
	s_in2(21,57)            <= s_out2(22,58);
	s_locks_lower_in(21,57) <= s_locks_lower_out(22,57);

		normal_cell_21_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,58),
			fetch              => s_fetch(21,58),
			data_in            => s_data_in(21,58),
			data_out           => s_data_out(21,58),
			out1               => s_out1(21,58),
			out2               => s_out2(21,58),
			lock_lower_row_out => s_locks_lower_out(21,58),
			lock_lower_row_in  => s_locks_lower_in(21,58),
			in1                => s_in1(21,58),
			in2                => s_in2(21,58),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(58)
		);
	s_in1(21,58)            <= s_out1(22,58);
	s_in2(21,58)            <= s_out2(22,59);
	s_locks_lower_in(21,58) <= s_locks_lower_out(22,58);

		normal_cell_21_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,59),
			fetch              => s_fetch(21,59),
			data_in            => s_data_in(21,59),
			data_out           => s_data_out(21,59),
			out1               => s_out1(21,59),
			out2               => s_out2(21,59),
			lock_lower_row_out => s_locks_lower_out(21,59),
			lock_lower_row_in  => s_locks_lower_in(21,59),
			in1                => s_in1(21,59),
			in2                => s_in2(21,59),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(59)
		);
	s_in1(21,59)            <= s_out1(22,59);
	s_in2(21,59)            <= s_out2(22,60);
	s_locks_lower_in(21,59) <= s_locks_lower_out(22,59);

		last_col_cell_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(21,60),
			fetch              => s_fetch(21,60),
			data_in            => s_data_in(21,60),
			data_out           => s_data_out(21,60),
			out1               => s_out1(21,60),
			out2               => s_out2(21,60),
			lock_lower_row_out => s_locks_lower_out(21,60),
			lock_lower_row_in  => s_locks_lower_in(21,60),
			in1                => s_in1(21,60),
			in2                => (others => '0'),
			lock_row           => s_locks(21),
			piv_found          => s_piv_found,
			row_data           => s_row_data(21),
			col_data           => s_col_data(60)
		);
	s_in1(21,60)            <= s_out1(22,60);
	s_locks_lower_in(21,60) <= s_locks_lower_out(22,60);

		normal_cell_22_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,1),
			fetch              => s_fetch(22,1),
			data_in            => s_data_in(22,1),
			data_out           => s_data_out(22,1),
			out1               => s_out1(22,1),
			out2               => s_out2(22,1),
			lock_lower_row_out => s_locks_lower_out(22,1),
			lock_lower_row_in  => s_locks_lower_in(22,1),
			in1                => s_in1(22,1),
			in2                => s_in2(22,1),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(1)
		);
	s_in1(22,1)            <= s_out1(23,1);
	s_in2(22,1)            <= s_out2(23,2);
	s_locks_lower_in(22,1) <= s_locks_lower_out(23,1);

		normal_cell_22_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,2),
			fetch              => s_fetch(22,2),
			data_in            => s_data_in(22,2),
			data_out           => s_data_out(22,2),
			out1               => s_out1(22,2),
			out2               => s_out2(22,2),
			lock_lower_row_out => s_locks_lower_out(22,2),
			lock_lower_row_in  => s_locks_lower_in(22,2),
			in1                => s_in1(22,2),
			in2                => s_in2(22,2),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(2)
		);
	s_in1(22,2)            <= s_out1(23,2);
	s_in2(22,2)            <= s_out2(23,3);
	s_locks_lower_in(22,2) <= s_locks_lower_out(23,2);

		normal_cell_22_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,3),
			fetch              => s_fetch(22,3),
			data_in            => s_data_in(22,3),
			data_out           => s_data_out(22,3),
			out1               => s_out1(22,3),
			out2               => s_out2(22,3),
			lock_lower_row_out => s_locks_lower_out(22,3),
			lock_lower_row_in  => s_locks_lower_in(22,3),
			in1                => s_in1(22,3),
			in2                => s_in2(22,3),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(3)
		);
	s_in1(22,3)            <= s_out1(23,3);
	s_in2(22,3)            <= s_out2(23,4);
	s_locks_lower_in(22,3) <= s_locks_lower_out(23,3);

		normal_cell_22_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,4),
			fetch              => s_fetch(22,4),
			data_in            => s_data_in(22,4),
			data_out           => s_data_out(22,4),
			out1               => s_out1(22,4),
			out2               => s_out2(22,4),
			lock_lower_row_out => s_locks_lower_out(22,4),
			lock_lower_row_in  => s_locks_lower_in(22,4),
			in1                => s_in1(22,4),
			in2                => s_in2(22,4),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(4)
		);
	s_in1(22,4)            <= s_out1(23,4);
	s_in2(22,4)            <= s_out2(23,5);
	s_locks_lower_in(22,4) <= s_locks_lower_out(23,4);

		normal_cell_22_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,5),
			fetch              => s_fetch(22,5),
			data_in            => s_data_in(22,5),
			data_out           => s_data_out(22,5),
			out1               => s_out1(22,5),
			out2               => s_out2(22,5),
			lock_lower_row_out => s_locks_lower_out(22,5),
			lock_lower_row_in  => s_locks_lower_in(22,5),
			in1                => s_in1(22,5),
			in2                => s_in2(22,5),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(5)
		);
	s_in1(22,5)            <= s_out1(23,5);
	s_in2(22,5)            <= s_out2(23,6);
	s_locks_lower_in(22,5) <= s_locks_lower_out(23,5);

		normal_cell_22_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,6),
			fetch              => s_fetch(22,6),
			data_in            => s_data_in(22,6),
			data_out           => s_data_out(22,6),
			out1               => s_out1(22,6),
			out2               => s_out2(22,6),
			lock_lower_row_out => s_locks_lower_out(22,6),
			lock_lower_row_in  => s_locks_lower_in(22,6),
			in1                => s_in1(22,6),
			in2                => s_in2(22,6),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(6)
		);
	s_in1(22,6)            <= s_out1(23,6);
	s_in2(22,6)            <= s_out2(23,7);
	s_locks_lower_in(22,6) <= s_locks_lower_out(23,6);

		normal_cell_22_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,7),
			fetch              => s_fetch(22,7),
			data_in            => s_data_in(22,7),
			data_out           => s_data_out(22,7),
			out1               => s_out1(22,7),
			out2               => s_out2(22,7),
			lock_lower_row_out => s_locks_lower_out(22,7),
			lock_lower_row_in  => s_locks_lower_in(22,7),
			in1                => s_in1(22,7),
			in2                => s_in2(22,7),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(7)
		);
	s_in1(22,7)            <= s_out1(23,7);
	s_in2(22,7)            <= s_out2(23,8);
	s_locks_lower_in(22,7) <= s_locks_lower_out(23,7);

		normal_cell_22_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,8),
			fetch              => s_fetch(22,8),
			data_in            => s_data_in(22,8),
			data_out           => s_data_out(22,8),
			out1               => s_out1(22,8),
			out2               => s_out2(22,8),
			lock_lower_row_out => s_locks_lower_out(22,8),
			lock_lower_row_in  => s_locks_lower_in(22,8),
			in1                => s_in1(22,8),
			in2                => s_in2(22,8),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(8)
		);
	s_in1(22,8)            <= s_out1(23,8);
	s_in2(22,8)            <= s_out2(23,9);
	s_locks_lower_in(22,8) <= s_locks_lower_out(23,8);

		normal_cell_22_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,9),
			fetch              => s_fetch(22,9),
			data_in            => s_data_in(22,9),
			data_out           => s_data_out(22,9),
			out1               => s_out1(22,9),
			out2               => s_out2(22,9),
			lock_lower_row_out => s_locks_lower_out(22,9),
			lock_lower_row_in  => s_locks_lower_in(22,9),
			in1                => s_in1(22,9),
			in2                => s_in2(22,9),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(9)
		);
	s_in1(22,9)            <= s_out1(23,9);
	s_in2(22,9)            <= s_out2(23,10);
	s_locks_lower_in(22,9) <= s_locks_lower_out(23,9);

		normal_cell_22_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,10),
			fetch              => s_fetch(22,10),
			data_in            => s_data_in(22,10),
			data_out           => s_data_out(22,10),
			out1               => s_out1(22,10),
			out2               => s_out2(22,10),
			lock_lower_row_out => s_locks_lower_out(22,10),
			lock_lower_row_in  => s_locks_lower_in(22,10),
			in1                => s_in1(22,10),
			in2                => s_in2(22,10),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(10)
		);
	s_in1(22,10)            <= s_out1(23,10);
	s_in2(22,10)            <= s_out2(23,11);
	s_locks_lower_in(22,10) <= s_locks_lower_out(23,10);

		normal_cell_22_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,11),
			fetch              => s_fetch(22,11),
			data_in            => s_data_in(22,11),
			data_out           => s_data_out(22,11),
			out1               => s_out1(22,11),
			out2               => s_out2(22,11),
			lock_lower_row_out => s_locks_lower_out(22,11),
			lock_lower_row_in  => s_locks_lower_in(22,11),
			in1                => s_in1(22,11),
			in2                => s_in2(22,11),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(11)
		);
	s_in1(22,11)            <= s_out1(23,11);
	s_in2(22,11)            <= s_out2(23,12);
	s_locks_lower_in(22,11) <= s_locks_lower_out(23,11);

		normal_cell_22_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,12),
			fetch              => s_fetch(22,12),
			data_in            => s_data_in(22,12),
			data_out           => s_data_out(22,12),
			out1               => s_out1(22,12),
			out2               => s_out2(22,12),
			lock_lower_row_out => s_locks_lower_out(22,12),
			lock_lower_row_in  => s_locks_lower_in(22,12),
			in1                => s_in1(22,12),
			in2                => s_in2(22,12),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(12)
		);
	s_in1(22,12)            <= s_out1(23,12);
	s_in2(22,12)            <= s_out2(23,13);
	s_locks_lower_in(22,12) <= s_locks_lower_out(23,12);

		normal_cell_22_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,13),
			fetch              => s_fetch(22,13),
			data_in            => s_data_in(22,13),
			data_out           => s_data_out(22,13),
			out1               => s_out1(22,13),
			out2               => s_out2(22,13),
			lock_lower_row_out => s_locks_lower_out(22,13),
			lock_lower_row_in  => s_locks_lower_in(22,13),
			in1                => s_in1(22,13),
			in2                => s_in2(22,13),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(13)
		);
	s_in1(22,13)            <= s_out1(23,13);
	s_in2(22,13)            <= s_out2(23,14);
	s_locks_lower_in(22,13) <= s_locks_lower_out(23,13);

		normal_cell_22_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,14),
			fetch              => s_fetch(22,14),
			data_in            => s_data_in(22,14),
			data_out           => s_data_out(22,14),
			out1               => s_out1(22,14),
			out2               => s_out2(22,14),
			lock_lower_row_out => s_locks_lower_out(22,14),
			lock_lower_row_in  => s_locks_lower_in(22,14),
			in1                => s_in1(22,14),
			in2                => s_in2(22,14),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(14)
		);
	s_in1(22,14)            <= s_out1(23,14);
	s_in2(22,14)            <= s_out2(23,15);
	s_locks_lower_in(22,14) <= s_locks_lower_out(23,14);

		normal_cell_22_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,15),
			fetch              => s_fetch(22,15),
			data_in            => s_data_in(22,15),
			data_out           => s_data_out(22,15),
			out1               => s_out1(22,15),
			out2               => s_out2(22,15),
			lock_lower_row_out => s_locks_lower_out(22,15),
			lock_lower_row_in  => s_locks_lower_in(22,15),
			in1                => s_in1(22,15),
			in2                => s_in2(22,15),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(15)
		);
	s_in1(22,15)            <= s_out1(23,15);
	s_in2(22,15)            <= s_out2(23,16);
	s_locks_lower_in(22,15) <= s_locks_lower_out(23,15);

		normal_cell_22_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,16),
			fetch              => s_fetch(22,16),
			data_in            => s_data_in(22,16),
			data_out           => s_data_out(22,16),
			out1               => s_out1(22,16),
			out2               => s_out2(22,16),
			lock_lower_row_out => s_locks_lower_out(22,16),
			lock_lower_row_in  => s_locks_lower_in(22,16),
			in1                => s_in1(22,16),
			in2                => s_in2(22,16),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(16)
		);
	s_in1(22,16)            <= s_out1(23,16);
	s_in2(22,16)            <= s_out2(23,17);
	s_locks_lower_in(22,16) <= s_locks_lower_out(23,16);

		normal_cell_22_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,17),
			fetch              => s_fetch(22,17),
			data_in            => s_data_in(22,17),
			data_out           => s_data_out(22,17),
			out1               => s_out1(22,17),
			out2               => s_out2(22,17),
			lock_lower_row_out => s_locks_lower_out(22,17),
			lock_lower_row_in  => s_locks_lower_in(22,17),
			in1                => s_in1(22,17),
			in2                => s_in2(22,17),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(17)
		);
	s_in1(22,17)            <= s_out1(23,17);
	s_in2(22,17)            <= s_out2(23,18);
	s_locks_lower_in(22,17) <= s_locks_lower_out(23,17);

		normal_cell_22_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,18),
			fetch              => s_fetch(22,18),
			data_in            => s_data_in(22,18),
			data_out           => s_data_out(22,18),
			out1               => s_out1(22,18),
			out2               => s_out2(22,18),
			lock_lower_row_out => s_locks_lower_out(22,18),
			lock_lower_row_in  => s_locks_lower_in(22,18),
			in1                => s_in1(22,18),
			in2                => s_in2(22,18),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(18)
		);
	s_in1(22,18)            <= s_out1(23,18);
	s_in2(22,18)            <= s_out2(23,19);
	s_locks_lower_in(22,18) <= s_locks_lower_out(23,18);

		normal_cell_22_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,19),
			fetch              => s_fetch(22,19),
			data_in            => s_data_in(22,19),
			data_out           => s_data_out(22,19),
			out1               => s_out1(22,19),
			out2               => s_out2(22,19),
			lock_lower_row_out => s_locks_lower_out(22,19),
			lock_lower_row_in  => s_locks_lower_in(22,19),
			in1                => s_in1(22,19),
			in2                => s_in2(22,19),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(19)
		);
	s_in1(22,19)            <= s_out1(23,19);
	s_in2(22,19)            <= s_out2(23,20);
	s_locks_lower_in(22,19) <= s_locks_lower_out(23,19);

		normal_cell_22_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,20),
			fetch              => s_fetch(22,20),
			data_in            => s_data_in(22,20),
			data_out           => s_data_out(22,20),
			out1               => s_out1(22,20),
			out2               => s_out2(22,20),
			lock_lower_row_out => s_locks_lower_out(22,20),
			lock_lower_row_in  => s_locks_lower_in(22,20),
			in1                => s_in1(22,20),
			in2                => s_in2(22,20),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(20)
		);
	s_in1(22,20)            <= s_out1(23,20);
	s_in2(22,20)            <= s_out2(23,21);
	s_locks_lower_in(22,20) <= s_locks_lower_out(23,20);

		normal_cell_22_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,21),
			fetch              => s_fetch(22,21),
			data_in            => s_data_in(22,21),
			data_out           => s_data_out(22,21),
			out1               => s_out1(22,21),
			out2               => s_out2(22,21),
			lock_lower_row_out => s_locks_lower_out(22,21),
			lock_lower_row_in  => s_locks_lower_in(22,21),
			in1                => s_in1(22,21),
			in2                => s_in2(22,21),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(21)
		);
	s_in1(22,21)            <= s_out1(23,21);
	s_in2(22,21)            <= s_out2(23,22);
	s_locks_lower_in(22,21) <= s_locks_lower_out(23,21);

		normal_cell_22_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,22),
			fetch              => s_fetch(22,22),
			data_in            => s_data_in(22,22),
			data_out           => s_data_out(22,22),
			out1               => s_out1(22,22),
			out2               => s_out2(22,22),
			lock_lower_row_out => s_locks_lower_out(22,22),
			lock_lower_row_in  => s_locks_lower_in(22,22),
			in1                => s_in1(22,22),
			in2                => s_in2(22,22),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(22)
		);
	s_in1(22,22)            <= s_out1(23,22);
	s_in2(22,22)            <= s_out2(23,23);
	s_locks_lower_in(22,22) <= s_locks_lower_out(23,22);

		normal_cell_22_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,23),
			fetch              => s_fetch(22,23),
			data_in            => s_data_in(22,23),
			data_out           => s_data_out(22,23),
			out1               => s_out1(22,23),
			out2               => s_out2(22,23),
			lock_lower_row_out => s_locks_lower_out(22,23),
			lock_lower_row_in  => s_locks_lower_in(22,23),
			in1                => s_in1(22,23),
			in2                => s_in2(22,23),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(23)
		);
	s_in1(22,23)            <= s_out1(23,23);
	s_in2(22,23)            <= s_out2(23,24);
	s_locks_lower_in(22,23) <= s_locks_lower_out(23,23);

		normal_cell_22_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,24),
			fetch              => s_fetch(22,24),
			data_in            => s_data_in(22,24),
			data_out           => s_data_out(22,24),
			out1               => s_out1(22,24),
			out2               => s_out2(22,24),
			lock_lower_row_out => s_locks_lower_out(22,24),
			lock_lower_row_in  => s_locks_lower_in(22,24),
			in1                => s_in1(22,24),
			in2                => s_in2(22,24),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(24)
		);
	s_in1(22,24)            <= s_out1(23,24);
	s_in2(22,24)            <= s_out2(23,25);
	s_locks_lower_in(22,24) <= s_locks_lower_out(23,24);

		normal_cell_22_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,25),
			fetch              => s_fetch(22,25),
			data_in            => s_data_in(22,25),
			data_out           => s_data_out(22,25),
			out1               => s_out1(22,25),
			out2               => s_out2(22,25),
			lock_lower_row_out => s_locks_lower_out(22,25),
			lock_lower_row_in  => s_locks_lower_in(22,25),
			in1                => s_in1(22,25),
			in2                => s_in2(22,25),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(25)
		);
	s_in1(22,25)            <= s_out1(23,25);
	s_in2(22,25)            <= s_out2(23,26);
	s_locks_lower_in(22,25) <= s_locks_lower_out(23,25);

		normal_cell_22_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,26),
			fetch              => s_fetch(22,26),
			data_in            => s_data_in(22,26),
			data_out           => s_data_out(22,26),
			out1               => s_out1(22,26),
			out2               => s_out2(22,26),
			lock_lower_row_out => s_locks_lower_out(22,26),
			lock_lower_row_in  => s_locks_lower_in(22,26),
			in1                => s_in1(22,26),
			in2                => s_in2(22,26),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(26)
		);
	s_in1(22,26)            <= s_out1(23,26);
	s_in2(22,26)            <= s_out2(23,27);
	s_locks_lower_in(22,26) <= s_locks_lower_out(23,26);

		normal_cell_22_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,27),
			fetch              => s_fetch(22,27),
			data_in            => s_data_in(22,27),
			data_out           => s_data_out(22,27),
			out1               => s_out1(22,27),
			out2               => s_out2(22,27),
			lock_lower_row_out => s_locks_lower_out(22,27),
			lock_lower_row_in  => s_locks_lower_in(22,27),
			in1                => s_in1(22,27),
			in2                => s_in2(22,27),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(27)
		);
	s_in1(22,27)            <= s_out1(23,27);
	s_in2(22,27)            <= s_out2(23,28);
	s_locks_lower_in(22,27) <= s_locks_lower_out(23,27);

		normal_cell_22_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,28),
			fetch              => s_fetch(22,28),
			data_in            => s_data_in(22,28),
			data_out           => s_data_out(22,28),
			out1               => s_out1(22,28),
			out2               => s_out2(22,28),
			lock_lower_row_out => s_locks_lower_out(22,28),
			lock_lower_row_in  => s_locks_lower_in(22,28),
			in1                => s_in1(22,28),
			in2                => s_in2(22,28),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(28)
		);
	s_in1(22,28)            <= s_out1(23,28);
	s_in2(22,28)            <= s_out2(23,29);
	s_locks_lower_in(22,28) <= s_locks_lower_out(23,28);

		normal_cell_22_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,29),
			fetch              => s_fetch(22,29),
			data_in            => s_data_in(22,29),
			data_out           => s_data_out(22,29),
			out1               => s_out1(22,29),
			out2               => s_out2(22,29),
			lock_lower_row_out => s_locks_lower_out(22,29),
			lock_lower_row_in  => s_locks_lower_in(22,29),
			in1                => s_in1(22,29),
			in2                => s_in2(22,29),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(29)
		);
	s_in1(22,29)            <= s_out1(23,29);
	s_in2(22,29)            <= s_out2(23,30);
	s_locks_lower_in(22,29) <= s_locks_lower_out(23,29);

		normal_cell_22_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,30),
			fetch              => s_fetch(22,30),
			data_in            => s_data_in(22,30),
			data_out           => s_data_out(22,30),
			out1               => s_out1(22,30),
			out2               => s_out2(22,30),
			lock_lower_row_out => s_locks_lower_out(22,30),
			lock_lower_row_in  => s_locks_lower_in(22,30),
			in1                => s_in1(22,30),
			in2                => s_in2(22,30),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(30)
		);
	s_in1(22,30)            <= s_out1(23,30);
	s_in2(22,30)            <= s_out2(23,31);
	s_locks_lower_in(22,30) <= s_locks_lower_out(23,30);

		normal_cell_22_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,31),
			fetch              => s_fetch(22,31),
			data_in            => s_data_in(22,31),
			data_out           => s_data_out(22,31),
			out1               => s_out1(22,31),
			out2               => s_out2(22,31),
			lock_lower_row_out => s_locks_lower_out(22,31),
			lock_lower_row_in  => s_locks_lower_in(22,31),
			in1                => s_in1(22,31),
			in2                => s_in2(22,31),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(31)
		);
	s_in1(22,31)            <= s_out1(23,31);
	s_in2(22,31)            <= s_out2(23,32);
	s_locks_lower_in(22,31) <= s_locks_lower_out(23,31);

		normal_cell_22_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,32),
			fetch              => s_fetch(22,32),
			data_in            => s_data_in(22,32),
			data_out           => s_data_out(22,32),
			out1               => s_out1(22,32),
			out2               => s_out2(22,32),
			lock_lower_row_out => s_locks_lower_out(22,32),
			lock_lower_row_in  => s_locks_lower_in(22,32),
			in1                => s_in1(22,32),
			in2                => s_in2(22,32),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(32)
		);
	s_in1(22,32)            <= s_out1(23,32);
	s_in2(22,32)            <= s_out2(23,33);
	s_locks_lower_in(22,32) <= s_locks_lower_out(23,32);

		normal_cell_22_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,33),
			fetch              => s_fetch(22,33),
			data_in            => s_data_in(22,33),
			data_out           => s_data_out(22,33),
			out1               => s_out1(22,33),
			out2               => s_out2(22,33),
			lock_lower_row_out => s_locks_lower_out(22,33),
			lock_lower_row_in  => s_locks_lower_in(22,33),
			in1                => s_in1(22,33),
			in2                => s_in2(22,33),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(33)
		);
	s_in1(22,33)            <= s_out1(23,33);
	s_in2(22,33)            <= s_out2(23,34);
	s_locks_lower_in(22,33) <= s_locks_lower_out(23,33);

		normal_cell_22_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,34),
			fetch              => s_fetch(22,34),
			data_in            => s_data_in(22,34),
			data_out           => s_data_out(22,34),
			out1               => s_out1(22,34),
			out2               => s_out2(22,34),
			lock_lower_row_out => s_locks_lower_out(22,34),
			lock_lower_row_in  => s_locks_lower_in(22,34),
			in1                => s_in1(22,34),
			in2                => s_in2(22,34),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(34)
		);
	s_in1(22,34)            <= s_out1(23,34);
	s_in2(22,34)            <= s_out2(23,35);
	s_locks_lower_in(22,34) <= s_locks_lower_out(23,34);

		normal_cell_22_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,35),
			fetch              => s_fetch(22,35),
			data_in            => s_data_in(22,35),
			data_out           => s_data_out(22,35),
			out1               => s_out1(22,35),
			out2               => s_out2(22,35),
			lock_lower_row_out => s_locks_lower_out(22,35),
			lock_lower_row_in  => s_locks_lower_in(22,35),
			in1                => s_in1(22,35),
			in2                => s_in2(22,35),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(35)
		);
	s_in1(22,35)            <= s_out1(23,35);
	s_in2(22,35)            <= s_out2(23,36);
	s_locks_lower_in(22,35) <= s_locks_lower_out(23,35);

		normal_cell_22_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,36),
			fetch              => s_fetch(22,36),
			data_in            => s_data_in(22,36),
			data_out           => s_data_out(22,36),
			out1               => s_out1(22,36),
			out2               => s_out2(22,36),
			lock_lower_row_out => s_locks_lower_out(22,36),
			lock_lower_row_in  => s_locks_lower_in(22,36),
			in1                => s_in1(22,36),
			in2                => s_in2(22,36),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(36)
		);
	s_in1(22,36)            <= s_out1(23,36);
	s_in2(22,36)            <= s_out2(23,37);
	s_locks_lower_in(22,36) <= s_locks_lower_out(23,36);

		normal_cell_22_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,37),
			fetch              => s_fetch(22,37),
			data_in            => s_data_in(22,37),
			data_out           => s_data_out(22,37),
			out1               => s_out1(22,37),
			out2               => s_out2(22,37),
			lock_lower_row_out => s_locks_lower_out(22,37),
			lock_lower_row_in  => s_locks_lower_in(22,37),
			in1                => s_in1(22,37),
			in2                => s_in2(22,37),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(37)
		);
	s_in1(22,37)            <= s_out1(23,37);
	s_in2(22,37)            <= s_out2(23,38);
	s_locks_lower_in(22,37) <= s_locks_lower_out(23,37);

		normal_cell_22_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,38),
			fetch              => s_fetch(22,38),
			data_in            => s_data_in(22,38),
			data_out           => s_data_out(22,38),
			out1               => s_out1(22,38),
			out2               => s_out2(22,38),
			lock_lower_row_out => s_locks_lower_out(22,38),
			lock_lower_row_in  => s_locks_lower_in(22,38),
			in1                => s_in1(22,38),
			in2                => s_in2(22,38),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(38)
		);
	s_in1(22,38)            <= s_out1(23,38);
	s_in2(22,38)            <= s_out2(23,39);
	s_locks_lower_in(22,38) <= s_locks_lower_out(23,38);

		normal_cell_22_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,39),
			fetch              => s_fetch(22,39),
			data_in            => s_data_in(22,39),
			data_out           => s_data_out(22,39),
			out1               => s_out1(22,39),
			out2               => s_out2(22,39),
			lock_lower_row_out => s_locks_lower_out(22,39),
			lock_lower_row_in  => s_locks_lower_in(22,39),
			in1                => s_in1(22,39),
			in2                => s_in2(22,39),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(39)
		);
	s_in1(22,39)            <= s_out1(23,39);
	s_in2(22,39)            <= s_out2(23,40);
	s_locks_lower_in(22,39) <= s_locks_lower_out(23,39);

		normal_cell_22_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,40),
			fetch              => s_fetch(22,40),
			data_in            => s_data_in(22,40),
			data_out           => s_data_out(22,40),
			out1               => s_out1(22,40),
			out2               => s_out2(22,40),
			lock_lower_row_out => s_locks_lower_out(22,40),
			lock_lower_row_in  => s_locks_lower_in(22,40),
			in1                => s_in1(22,40),
			in2                => s_in2(22,40),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(40)
		);
	s_in1(22,40)            <= s_out1(23,40);
	s_in2(22,40)            <= s_out2(23,41);
	s_locks_lower_in(22,40) <= s_locks_lower_out(23,40);

		normal_cell_22_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,41),
			fetch              => s_fetch(22,41),
			data_in            => s_data_in(22,41),
			data_out           => s_data_out(22,41),
			out1               => s_out1(22,41),
			out2               => s_out2(22,41),
			lock_lower_row_out => s_locks_lower_out(22,41),
			lock_lower_row_in  => s_locks_lower_in(22,41),
			in1                => s_in1(22,41),
			in2                => s_in2(22,41),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(41)
		);
	s_in1(22,41)            <= s_out1(23,41);
	s_in2(22,41)            <= s_out2(23,42);
	s_locks_lower_in(22,41) <= s_locks_lower_out(23,41);

		normal_cell_22_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,42),
			fetch              => s_fetch(22,42),
			data_in            => s_data_in(22,42),
			data_out           => s_data_out(22,42),
			out1               => s_out1(22,42),
			out2               => s_out2(22,42),
			lock_lower_row_out => s_locks_lower_out(22,42),
			lock_lower_row_in  => s_locks_lower_in(22,42),
			in1                => s_in1(22,42),
			in2                => s_in2(22,42),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(42)
		);
	s_in1(22,42)            <= s_out1(23,42);
	s_in2(22,42)            <= s_out2(23,43);
	s_locks_lower_in(22,42) <= s_locks_lower_out(23,42);

		normal_cell_22_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,43),
			fetch              => s_fetch(22,43),
			data_in            => s_data_in(22,43),
			data_out           => s_data_out(22,43),
			out1               => s_out1(22,43),
			out2               => s_out2(22,43),
			lock_lower_row_out => s_locks_lower_out(22,43),
			lock_lower_row_in  => s_locks_lower_in(22,43),
			in1                => s_in1(22,43),
			in2                => s_in2(22,43),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(43)
		);
	s_in1(22,43)            <= s_out1(23,43);
	s_in2(22,43)            <= s_out2(23,44);
	s_locks_lower_in(22,43) <= s_locks_lower_out(23,43);

		normal_cell_22_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,44),
			fetch              => s_fetch(22,44),
			data_in            => s_data_in(22,44),
			data_out           => s_data_out(22,44),
			out1               => s_out1(22,44),
			out2               => s_out2(22,44),
			lock_lower_row_out => s_locks_lower_out(22,44),
			lock_lower_row_in  => s_locks_lower_in(22,44),
			in1                => s_in1(22,44),
			in2                => s_in2(22,44),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(44)
		);
	s_in1(22,44)            <= s_out1(23,44);
	s_in2(22,44)            <= s_out2(23,45);
	s_locks_lower_in(22,44) <= s_locks_lower_out(23,44);

		normal_cell_22_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,45),
			fetch              => s_fetch(22,45),
			data_in            => s_data_in(22,45),
			data_out           => s_data_out(22,45),
			out1               => s_out1(22,45),
			out2               => s_out2(22,45),
			lock_lower_row_out => s_locks_lower_out(22,45),
			lock_lower_row_in  => s_locks_lower_in(22,45),
			in1                => s_in1(22,45),
			in2                => s_in2(22,45),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(45)
		);
	s_in1(22,45)            <= s_out1(23,45);
	s_in2(22,45)            <= s_out2(23,46);
	s_locks_lower_in(22,45) <= s_locks_lower_out(23,45);

		normal_cell_22_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,46),
			fetch              => s_fetch(22,46),
			data_in            => s_data_in(22,46),
			data_out           => s_data_out(22,46),
			out1               => s_out1(22,46),
			out2               => s_out2(22,46),
			lock_lower_row_out => s_locks_lower_out(22,46),
			lock_lower_row_in  => s_locks_lower_in(22,46),
			in1                => s_in1(22,46),
			in2                => s_in2(22,46),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(46)
		);
	s_in1(22,46)            <= s_out1(23,46);
	s_in2(22,46)            <= s_out2(23,47);
	s_locks_lower_in(22,46) <= s_locks_lower_out(23,46);

		normal_cell_22_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,47),
			fetch              => s_fetch(22,47),
			data_in            => s_data_in(22,47),
			data_out           => s_data_out(22,47),
			out1               => s_out1(22,47),
			out2               => s_out2(22,47),
			lock_lower_row_out => s_locks_lower_out(22,47),
			lock_lower_row_in  => s_locks_lower_in(22,47),
			in1                => s_in1(22,47),
			in2                => s_in2(22,47),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(47)
		);
	s_in1(22,47)            <= s_out1(23,47);
	s_in2(22,47)            <= s_out2(23,48);
	s_locks_lower_in(22,47) <= s_locks_lower_out(23,47);

		normal_cell_22_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,48),
			fetch              => s_fetch(22,48),
			data_in            => s_data_in(22,48),
			data_out           => s_data_out(22,48),
			out1               => s_out1(22,48),
			out2               => s_out2(22,48),
			lock_lower_row_out => s_locks_lower_out(22,48),
			lock_lower_row_in  => s_locks_lower_in(22,48),
			in1                => s_in1(22,48),
			in2                => s_in2(22,48),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(48)
		);
	s_in1(22,48)            <= s_out1(23,48);
	s_in2(22,48)            <= s_out2(23,49);
	s_locks_lower_in(22,48) <= s_locks_lower_out(23,48);

		normal_cell_22_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,49),
			fetch              => s_fetch(22,49),
			data_in            => s_data_in(22,49),
			data_out           => s_data_out(22,49),
			out1               => s_out1(22,49),
			out2               => s_out2(22,49),
			lock_lower_row_out => s_locks_lower_out(22,49),
			lock_lower_row_in  => s_locks_lower_in(22,49),
			in1                => s_in1(22,49),
			in2                => s_in2(22,49),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(49)
		);
	s_in1(22,49)            <= s_out1(23,49);
	s_in2(22,49)            <= s_out2(23,50);
	s_locks_lower_in(22,49) <= s_locks_lower_out(23,49);

		normal_cell_22_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,50),
			fetch              => s_fetch(22,50),
			data_in            => s_data_in(22,50),
			data_out           => s_data_out(22,50),
			out1               => s_out1(22,50),
			out2               => s_out2(22,50),
			lock_lower_row_out => s_locks_lower_out(22,50),
			lock_lower_row_in  => s_locks_lower_in(22,50),
			in1                => s_in1(22,50),
			in2                => s_in2(22,50),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(50)
		);
	s_in1(22,50)            <= s_out1(23,50);
	s_in2(22,50)            <= s_out2(23,51);
	s_locks_lower_in(22,50) <= s_locks_lower_out(23,50);

		normal_cell_22_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,51),
			fetch              => s_fetch(22,51),
			data_in            => s_data_in(22,51),
			data_out           => s_data_out(22,51),
			out1               => s_out1(22,51),
			out2               => s_out2(22,51),
			lock_lower_row_out => s_locks_lower_out(22,51),
			lock_lower_row_in  => s_locks_lower_in(22,51),
			in1                => s_in1(22,51),
			in2                => s_in2(22,51),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(51)
		);
	s_in1(22,51)            <= s_out1(23,51);
	s_in2(22,51)            <= s_out2(23,52);
	s_locks_lower_in(22,51) <= s_locks_lower_out(23,51);

		normal_cell_22_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,52),
			fetch              => s_fetch(22,52),
			data_in            => s_data_in(22,52),
			data_out           => s_data_out(22,52),
			out1               => s_out1(22,52),
			out2               => s_out2(22,52),
			lock_lower_row_out => s_locks_lower_out(22,52),
			lock_lower_row_in  => s_locks_lower_in(22,52),
			in1                => s_in1(22,52),
			in2                => s_in2(22,52),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(52)
		);
	s_in1(22,52)            <= s_out1(23,52);
	s_in2(22,52)            <= s_out2(23,53);
	s_locks_lower_in(22,52) <= s_locks_lower_out(23,52);

		normal_cell_22_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,53),
			fetch              => s_fetch(22,53),
			data_in            => s_data_in(22,53),
			data_out           => s_data_out(22,53),
			out1               => s_out1(22,53),
			out2               => s_out2(22,53),
			lock_lower_row_out => s_locks_lower_out(22,53),
			lock_lower_row_in  => s_locks_lower_in(22,53),
			in1                => s_in1(22,53),
			in2                => s_in2(22,53),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(53)
		);
	s_in1(22,53)            <= s_out1(23,53);
	s_in2(22,53)            <= s_out2(23,54);
	s_locks_lower_in(22,53) <= s_locks_lower_out(23,53);

		normal_cell_22_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,54),
			fetch              => s_fetch(22,54),
			data_in            => s_data_in(22,54),
			data_out           => s_data_out(22,54),
			out1               => s_out1(22,54),
			out2               => s_out2(22,54),
			lock_lower_row_out => s_locks_lower_out(22,54),
			lock_lower_row_in  => s_locks_lower_in(22,54),
			in1                => s_in1(22,54),
			in2                => s_in2(22,54),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(54)
		);
	s_in1(22,54)            <= s_out1(23,54);
	s_in2(22,54)            <= s_out2(23,55);
	s_locks_lower_in(22,54) <= s_locks_lower_out(23,54);

		normal_cell_22_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,55),
			fetch              => s_fetch(22,55),
			data_in            => s_data_in(22,55),
			data_out           => s_data_out(22,55),
			out1               => s_out1(22,55),
			out2               => s_out2(22,55),
			lock_lower_row_out => s_locks_lower_out(22,55),
			lock_lower_row_in  => s_locks_lower_in(22,55),
			in1                => s_in1(22,55),
			in2                => s_in2(22,55),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(55)
		);
	s_in1(22,55)            <= s_out1(23,55);
	s_in2(22,55)            <= s_out2(23,56);
	s_locks_lower_in(22,55) <= s_locks_lower_out(23,55);

		normal_cell_22_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,56),
			fetch              => s_fetch(22,56),
			data_in            => s_data_in(22,56),
			data_out           => s_data_out(22,56),
			out1               => s_out1(22,56),
			out2               => s_out2(22,56),
			lock_lower_row_out => s_locks_lower_out(22,56),
			lock_lower_row_in  => s_locks_lower_in(22,56),
			in1                => s_in1(22,56),
			in2                => s_in2(22,56),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(56)
		);
	s_in1(22,56)            <= s_out1(23,56);
	s_in2(22,56)            <= s_out2(23,57);
	s_locks_lower_in(22,56) <= s_locks_lower_out(23,56);

		normal_cell_22_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,57),
			fetch              => s_fetch(22,57),
			data_in            => s_data_in(22,57),
			data_out           => s_data_out(22,57),
			out1               => s_out1(22,57),
			out2               => s_out2(22,57),
			lock_lower_row_out => s_locks_lower_out(22,57),
			lock_lower_row_in  => s_locks_lower_in(22,57),
			in1                => s_in1(22,57),
			in2                => s_in2(22,57),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(57)
		);
	s_in1(22,57)            <= s_out1(23,57);
	s_in2(22,57)            <= s_out2(23,58);
	s_locks_lower_in(22,57) <= s_locks_lower_out(23,57);

		normal_cell_22_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,58),
			fetch              => s_fetch(22,58),
			data_in            => s_data_in(22,58),
			data_out           => s_data_out(22,58),
			out1               => s_out1(22,58),
			out2               => s_out2(22,58),
			lock_lower_row_out => s_locks_lower_out(22,58),
			lock_lower_row_in  => s_locks_lower_in(22,58),
			in1                => s_in1(22,58),
			in2                => s_in2(22,58),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(58)
		);
	s_in1(22,58)            <= s_out1(23,58);
	s_in2(22,58)            <= s_out2(23,59);
	s_locks_lower_in(22,58) <= s_locks_lower_out(23,58);

		normal_cell_22_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,59),
			fetch              => s_fetch(22,59),
			data_in            => s_data_in(22,59),
			data_out           => s_data_out(22,59),
			out1               => s_out1(22,59),
			out2               => s_out2(22,59),
			lock_lower_row_out => s_locks_lower_out(22,59),
			lock_lower_row_in  => s_locks_lower_in(22,59),
			in1                => s_in1(22,59),
			in2                => s_in2(22,59),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(59)
		);
	s_in1(22,59)            <= s_out1(23,59);
	s_in2(22,59)            <= s_out2(23,60);
	s_locks_lower_in(22,59) <= s_locks_lower_out(23,59);

		last_col_cell_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(22,60),
			fetch              => s_fetch(22,60),
			data_in            => s_data_in(22,60),
			data_out           => s_data_out(22,60),
			out1               => s_out1(22,60),
			out2               => s_out2(22,60),
			lock_lower_row_out => s_locks_lower_out(22,60),
			lock_lower_row_in  => s_locks_lower_in(22,60),
			in1                => s_in1(22,60),
			in2                => (others => '0'),
			lock_row           => s_locks(22),
			piv_found          => s_piv_found,
			row_data           => s_row_data(22),
			col_data           => s_col_data(60)
		);
	s_in1(22,60)            <= s_out1(23,60);
	s_locks_lower_in(22,60) <= s_locks_lower_out(23,60);

		normal_cell_23_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,1),
			fetch              => s_fetch(23,1),
			data_in            => s_data_in(23,1),
			data_out           => s_data_out(23,1),
			out1               => s_out1(23,1),
			out2               => s_out2(23,1),
			lock_lower_row_out => s_locks_lower_out(23,1),
			lock_lower_row_in  => s_locks_lower_in(23,1),
			in1                => s_in1(23,1),
			in2                => s_in2(23,1),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(1)
		);
	s_in1(23,1)            <= s_out1(24,1);
	s_in2(23,1)            <= s_out2(24,2);
	s_locks_lower_in(23,1) <= s_locks_lower_out(24,1);

		normal_cell_23_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,2),
			fetch              => s_fetch(23,2),
			data_in            => s_data_in(23,2),
			data_out           => s_data_out(23,2),
			out1               => s_out1(23,2),
			out2               => s_out2(23,2),
			lock_lower_row_out => s_locks_lower_out(23,2),
			lock_lower_row_in  => s_locks_lower_in(23,2),
			in1                => s_in1(23,2),
			in2                => s_in2(23,2),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(2)
		);
	s_in1(23,2)            <= s_out1(24,2);
	s_in2(23,2)            <= s_out2(24,3);
	s_locks_lower_in(23,2) <= s_locks_lower_out(24,2);

		normal_cell_23_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,3),
			fetch              => s_fetch(23,3),
			data_in            => s_data_in(23,3),
			data_out           => s_data_out(23,3),
			out1               => s_out1(23,3),
			out2               => s_out2(23,3),
			lock_lower_row_out => s_locks_lower_out(23,3),
			lock_lower_row_in  => s_locks_lower_in(23,3),
			in1                => s_in1(23,3),
			in2                => s_in2(23,3),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(3)
		);
	s_in1(23,3)            <= s_out1(24,3);
	s_in2(23,3)            <= s_out2(24,4);
	s_locks_lower_in(23,3) <= s_locks_lower_out(24,3);

		normal_cell_23_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,4),
			fetch              => s_fetch(23,4),
			data_in            => s_data_in(23,4),
			data_out           => s_data_out(23,4),
			out1               => s_out1(23,4),
			out2               => s_out2(23,4),
			lock_lower_row_out => s_locks_lower_out(23,4),
			lock_lower_row_in  => s_locks_lower_in(23,4),
			in1                => s_in1(23,4),
			in2                => s_in2(23,4),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(4)
		);
	s_in1(23,4)            <= s_out1(24,4);
	s_in2(23,4)            <= s_out2(24,5);
	s_locks_lower_in(23,4) <= s_locks_lower_out(24,4);

		normal_cell_23_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,5),
			fetch              => s_fetch(23,5),
			data_in            => s_data_in(23,5),
			data_out           => s_data_out(23,5),
			out1               => s_out1(23,5),
			out2               => s_out2(23,5),
			lock_lower_row_out => s_locks_lower_out(23,5),
			lock_lower_row_in  => s_locks_lower_in(23,5),
			in1                => s_in1(23,5),
			in2                => s_in2(23,5),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(5)
		);
	s_in1(23,5)            <= s_out1(24,5);
	s_in2(23,5)            <= s_out2(24,6);
	s_locks_lower_in(23,5) <= s_locks_lower_out(24,5);

		normal_cell_23_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,6),
			fetch              => s_fetch(23,6),
			data_in            => s_data_in(23,6),
			data_out           => s_data_out(23,6),
			out1               => s_out1(23,6),
			out2               => s_out2(23,6),
			lock_lower_row_out => s_locks_lower_out(23,6),
			lock_lower_row_in  => s_locks_lower_in(23,6),
			in1                => s_in1(23,6),
			in2                => s_in2(23,6),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(6)
		);
	s_in1(23,6)            <= s_out1(24,6);
	s_in2(23,6)            <= s_out2(24,7);
	s_locks_lower_in(23,6) <= s_locks_lower_out(24,6);

		normal_cell_23_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,7),
			fetch              => s_fetch(23,7),
			data_in            => s_data_in(23,7),
			data_out           => s_data_out(23,7),
			out1               => s_out1(23,7),
			out2               => s_out2(23,7),
			lock_lower_row_out => s_locks_lower_out(23,7),
			lock_lower_row_in  => s_locks_lower_in(23,7),
			in1                => s_in1(23,7),
			in2                => s_in2(23,7),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(7)
		);
	s_in1(23,7)            <= s_out1(24,7);
	s_in2(23,7)            <= s_out2(24,8);
	s_locks_lower_in(23,7) <= s_locks_lower_out(24,7);

		normal_cell_23_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,8),
			fetch              => s_fetch(23,8),
			data_in            => s_data_in(23,8),
			data_out           => s_data_out(23,8),
			out1               => s_out1(23,8),
			out2               => s_out2(23,8),
			lock_lower_row_out => s_locks_lower_out(23,8),
			lock_lower_row_in  => s_locks_lower_in(23,8),
			in1                => s_in1(23,8),
			in2                => s_in2(23,8),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(8)
		);
	s_in1(23,8)            <= s_out1(24,8);
	s_in2(23,8)            <= s_out2(24,9);
	s_locks_lower_in(23,8) <= s_locks_lower_out(24,8);

		normal_cell_23_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,9),
			fetch              => s_fetch(23,9),
			data_in            => s_data_in(23,9),
			data_out           => s_data_out(23,9),
			out1               => s_out1(23,9),
			out2               => s_out2(23,9),
			lock_lower_row_out => s_locks_lower_out(23,9),
			lock_lower_row_in  => s_locks_lower_in(23,9),
			in1                => s_in1(23,9),
			in2                => s_in2(23,9),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(9)
		);
	s_in1(23,9)            <= s_out1(24,9);
	s_in2(23,9)            <= s_out2(24,10);
	s_locks_lower_in(23,9) <= s_locks_lower_out(24,9);

		normal_cell_23_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,10),
			fetch              => s_fetch(23,10),
			data_in            => s_data_in(23,10),
			data_out           => s_data_out(23,10),
			out1               => s_out1(23,10),
			out2               => s_out2(23,10),
			lock_lower_row_out => s_locks_lower_out(23,10),
			lock_lower_row_in  => s_locks_lower_in(23,10),
			in1                => s_in1(23,10),
			in2                => s_in2(23,10),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(10)
		);
	s_in1(23,10)            <= s_out1(24,10);
	s_in2(23,10)            <= s_out2(24,11);
	s_locks_lower_in(23,10) <= s_locks_lower_out(24,10);

		normal_cell_23_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,11),
			fetch              => s_fetch(23,11),
			data_in            => s_data_in(23,11),
			data_out           => s_data_out(23,11),
			out1               => s_out1(23,11),
			out2               => s_out2(23,11),
			lock_lower_row_out => s_locks_lower_out(23,11),
			lock_lower_row_in  => s_locks_lower_in(23,11),
			in1                => s_in1(23,11),
			in2                => s_in2(23,11),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(11)
		);
	s_in1(23,11)            <= s_out1(24,11);
	s_in2(23,11)            <= s_out2(24,12);
	s_locks_lower_in(23,11) <= s_locks_lower_out(24,11);

		normal_cell_23_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,12),
			fetch              => s_fetch(23,12),
			data_in            => s_data_in(23,12),
			data_out           => s_data_out(23,12),
			out1               => s_out1(23,12),
			out2               => s_out2(23,12),
			lock_lower_row_out => s_locks_lower_out(23,12),
			lock_lower_row_in  => s_locks_lower_in(23,12),
			in1                => s_in1(23,12),
			in2                => s_in2(23,12),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(12)
		);
	s_in1(23,12)            <= s_out1(24,12);
	s_in2(23,12)            <= s_out2(24,13);
	s_locks_lower_in(23,12) <= s_locks_lower_out(24,12);

		normal_cell_23_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,13),
			fetch              => s_fetch(23,13),
			data_in            => s_data_in(23,13),
			data_out           => s_data_out(23,13),
			out1               => s_out1(23,13),
			out2               => s_out2(23,13),
			lock_lower_row_out => s_locks_lower_out(23,13),
			lock_lower_row_in  => s_locks_lower_in(23,13),
			in1                => s_in1(23,13),
			in2                => s_in2(23,13),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(13)
		);
	s_in1(23,13)            <= s_out1(24,13);
	s_in2(23,13)            <= s_out2(24,14);
	s_locks_lower_in(23,13) <= s_locks_lower_out(24,13);

		normal_cell_23_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,14),
			fetch              => s_fetch(23,14),
			data_in            => s_data_in(23,14),
			data_out           => s_data_out(23,14),
			out1               => s_out1(23,14),
			out2               => s_out2(23,14),
			lock_lower_row_out => s_locks_lower_out(23,14),
			lock_lower_row_in  => s_locks_lower_in(23,14),
			in1                => s_in1(23,14),
			in2                => s_in2(23,14),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(14)
		);
	s_in1(23,14)            <= s_out1(24,14);
	s_in2(23,14)            <= s_out2(24,15);
	s_locks_lower_in(23,14) <= s_locks_lower_out(24,14);

		normal_cell_23_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,15),
			fetch              => s_fetch(23,15),
			data_in            => s_data_in(23,15),
			data_out           => s_data_out(23,15),
			out1               => s_out1(23,15),
			out2               => s_out2(23,15),
			lock_lower_row_out => s_locks_lower_out(23,15),
			lock_lower_row_in  => s_locks_lower_in(23,15),
			in1                => s_in1(23,15),
			in2                => s_in2(23,15),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(15)
		);
	s_in1(23,15)            <= s_out1(24,15);
	s_in2(23,15)            <= s_out2(24,16);
	s_locks_lower_in(23,15) <= s_locks_lower_out(24,15);

		normal_cell_23_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,16),
			fetch              => s_fetch(23,16),
			data_in            => s_data_in(23,16),
			data_out           => s_data_out(23,16),
			out1               => s_out1(23,16),
			out2               => s_out2(23,16),
			lock_lower_row_out => s_locks_lower_out(23,16),
			lock_lower_row_in  => s_locks_lower_in(23,16),
			in1                => s_in1(23,16),
			in2                => s_in2(23,16),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(16)
		);
	s_in1(23,16)            <= s_out1(24,16);
	s_in2(23,16)            <= s_out2(24,17);
	s_locks_lower_in(23,16) <= s_locks_lower_out(24,16);

		normal_cell_23_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,17),
			fetch              => s_fetch(23,17),
			data_in            => s_data_in(23,17),
			data_out           => s_data_out(23,17),
			out1               => s_out1(23,17),
			out2               => s_out2(23,17),
			lock_lower_row_out => s_locks_lower_out(23,17),
			lock_lower_row_in  => s_locks_lower_in(23,17),
			in1                => s_in1(23,17),
			in2                => s_in2(23,17),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(17)
		);
	s_in1(23,17)            <= s_out1(24,17);
	s_in2(23,17)            <= s_out2(24,18);
	s_locks_lower_in(23,17) <= s_locks_lower_out(24,17);

		normal_cell_23_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,18),
			fetch              => s_fetch(23,18),
			data_in            => s_data_in(23,18),
			data_out           => s_data_out(23,18),
			out1               => s_out1(23,18),
			out2               => s_out2(23,18),
			lock_lower_row_out => s_locks_lower_out(23,18),
			lock_lower_row_in  => s_locks_lower_in(23,18),
			in1                => s_in1(23,18),
			in2                => s_in2(23,18),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(18)
		);
	s_in1(23,18)            <= s_out1(24,18);
	s_in2(23,18)            <= s_out2(24,19);
	s_locks_lower_in(23,18) <= s_locks_lower_out(24,18);

		normal_cell_23_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,19),
			fetch              => s_fetch(23,19),
			data_in            => s_data_in(23,19),
			data_out           => s_data_out(23,19),
			out1               => s_out1(23,19),
			out2               => s_out2(23,19),
			lock_lower_row_out => s_locks_lower_out(23,19),
			lock_lower_row_in  => s_locks_lower_in(23,19),
			in1                => s_in1(23,19),
			in2                => s_in2(23,19),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(19)
		);
	s_in1(23,19)            <= s_out1(24,19);
	s_in2(23,19)            <= s_out2(24,20);
	s_locks_lower_in(23,19) <= s_locks_lower_out(24,19);

		normal_cell_23_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,20),
			fetch              => s_fetch(23,20),
			data_in            => s_data_in(23,20),
			data_out           => s_data_out(23,20),
			out1               => s_out1(23,20),
			out2               => s_out2(23,20),
			lock_lower_row_out => s_locks_lower_out(23,20),
			lock_lower_row_in  => s_locks_lower_in(23,20),
			in1                => s_in1(23,20),
			in2                => s_in2(23,20),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(20)
		);
	s_in1(23,20)            <= s_out1(24,20);
	s_in2(23,20)            <= s_out2(24,21);
	s_locks_lower_in(23,20) <= s_locks_lower_out(24,20);

		normal_cell_23_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,21),
			fetch              => s_fetch(23,21),
			data_in            => s_data_in(23,21),
			data_out           => s_data_out(23,21),
			out1               => s_out1(23,21),
			out2               => s_out2(23,21),
			lock_lower_row_out => s_locks_lower_out(23,21),
			lock_lower_row_in  => s_locks_lower_in(23,21),
			in1                => s_in1(23,21),
			in2                => s_in2(23,21),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(21)
		);
	s_in1(23,21)            <= s_out1(24,21);
	s_in2(23,21)            <= s_out2(24,22);
	s_locks_lower_in(23,21) <= s_locks_lower_out(24,21);

		normal_cell_23_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,22),
			fetch              => s_fetch(23,22),
			data_in            => s_data_in(23,22),
			data_out           => s_data_out(23,22),
			out1               => s_out1(23,22),
			out2               => s_out2(23,22),
			lock_lower_row_out => s_locks_lower_out(23,22),
			lock_lower_row_in  => s_locks_lower_in(23,22),
			in1                => s_in1(23,22),
			in2                => s_in2(23,22),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(22)
		);
	s_in1(23,22)            <= s_out1(24,22);
	s_in2(23,22)            <= s_out2(24,23);
	s_locks_lower_in(23,22) <= s_locks_lower_out(24,22);

		normal_cell_23_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,23),
			fetch              => s_fetch(23,23),
			data_in            => s_data_in(23,23),
			data_out           => s_data_out(23,23),
			out1               => s_out1(23,23),
			out2               => s_out2(23,23),
			lock_lower_row_out => s_locks_lower_out(23,23),
			lock_lower_row_in  => s_locks_lower_in(23,23),
			in1                => s_in1(23,23),
			in2                => s_in2(23,23),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(23)
		);
	s_in1(23,23)            <= s_out1(24,23);
	s_in2(23,23)            <= s_out2(24,24);
	s_locks_lower_in(23,23) <= s_locks_lower_out(24,23);

		normal_cell_23_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,24),
			fetch              => s_fetch(23,24),
			data_in            => s_data_in(23,24),
			data_out           => s_data_out(23,24),
			out1               => s_out1(23,24),
			out2               => s_out2(23,24),
			lock_lower_row_out => s_locks_lower_out(23,24),
			lock_lower_row_in  => s_locks_lower_in(23,24),
			in1                => s_in1(23,24),
			in2                => s_in2(23,24),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(24)
		);
	s_in1(23,24)            <= s_out1(24,24);
	s_in2(23,24)            <= s_out2(24,25);
	s_locks_lower_in(23,24) <= s_locks_lower_out(24,24);

		normal_cell_23_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,25),
			fetch              => s_fetch(23,25),
			data_in            => s_data_in(23,25),
			data_out           => s_data_out(23,25),
			out1               => s_out1(23,25),
			out2               => s_out2(23,25),
			lock_lower_row_out => s_locks_lower_out(23,25),
			lock_lower_row_in  => s_locks_lower_in(23,25),
			in1                => s_in1(23,25),
			in2                => s_in2(23,25),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(25)
		);
	s_in1(23,25)            <= s_out1(24,25);
	s_in2(23,25)            <= s_out2(24,26);
	s_locks_lower_in(23,25) <= s_locks_lower_out(24,25);

		normal_cell_23_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,26),
			fetch              => s_fetch(23,26),
			data_in            => s_data_in(23,26),
			data_out           => s_data_out(23,26),
			out1               => s_out1(23,26),
			out2               => s_out2(23,26),
			lock_lower_row_out => s_locks_lower_out(23,26),
			lock_lower_row_in  => s_locks_lower_in(23,26),
			in1                => s_in1(23,26),
			in2                => s_in2(23,26),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(26)
		);
	s_in1(23,26)            <= s_out1(24,26);
	s_in2(23,26)            <= s_out2(24,27);
	s_locks_lower_in(23,26) <= s_locks_lower_out(24,26);

		normal_cell_23_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,27),
			fetch              => s_fetch(23,27),
			data_in            => s_data_in(23,27),
			data_out           => s_data_out(23,27),
			out1               => s_out1(23,27),
			out2               => s_out2(23,27),
			lock_lower_row_out => s_locks_lower_out(23,27),
			lock_lower_row_in  => s_locks_lower_in(23,27),
			in1                => s_in1(23,27),
			in2                => s_in2(23,27),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(27)
		);
	s_in1(23,27)            <= s_out1(24,27);
	s_in2(23,27)            <= s_out2(24,28);
	s_locks_lower_in(23,27) <= s_locks_lower_out(24,27);

		normal_cell_23_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,28),
			fetch              => s_fetch(23,28),
			data_in            => s_data_in(23,28),
			data_out           => s_data_out(23,28),
			out1               => s_out1(23,28),
			out2               => s_out2(23,28),
			lock_lower_row_out => s_locks_lower_out(23,28),
			lock_lower_row_in  => s_locks_lower_in(23,28),
			in1                => s_in1(23,28),
			in2                => s_in2(23,28),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(28)
		);
	s_in1(23,28)            <= s_out1(24,28);
	s_in2(23,28)            <= s_out2(24,29);
	s_locks_lower_in(23,28) <= s_locks_lower_out(24,28);

		normal_cell_23_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,29),
			fetch              => s_fetch(23,29),
			data_in            => s_data_in(23,29),
			data_out           => s_data_out(23,29),
			out1               => s_out1(23,29),
			out2               => s_out2(23,29),
			lock_lower_row_out => s_locks_lower_out(23,29),
			lock_lower_row_in  => s_locks_lower_in(23,29),
			in1                => s_in1(23,29),
			in2                => s_in2(23,29),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(29)
		);
	s_in1(23,29)            <= s_out1(24,29);
	s_in2(23,29)            <= s_out2(24,30);
	s_locks_lower_in(23,29) <= s_locks_lower_out(24,29);

		normal_cell_23_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,30),
			fetch              => s_fetch(23,30),
			data_in            => s_data_in(23,30),
			data_out           => s_data_out(23,30),
			out1               => s_out1(23,30),
			out2               => s_out2(23,30),
			lock_lower_row_out => s_locks_lower_out(23,30),
			lock_lower_row_in  => s_locks_lower_in(23,30),
			in1                => s_in1(23,30),
			in2                => s_in2(23,30),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(30)
		);
	s_in1(23,30)            <= s_out1(24,30);
	s_in2(23,30)            <= s_out2(24,31);
	s_locks_lower_in(23,30) <= s_locks_lower_out(24,30);

		normal_cell_23_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,31),
			fetch              => s_fetch(23,31),
			data_in            => s_data_in(23,31),
			data_out           => s_data_out(23,31),
			out1               => s_out1(23,31),
			out2               => s_out2(23,31),
			lock_lower_row_out => s_locks_lower_out(23,31),
			lock_lower_row_in  => s_locks_lower_in(23,31),
			in1                => s_in1(23,31),
			in2                => s_in2(23,31),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(31)
		);
	s_in1(23,31)            <= s_out1(24,31);
	s_in2(23,31)            <= s_out2(24,32);
	s_locks_lower_in(23,31) <= s_locks_lower_out(24,31);

		normal_cell_23_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,32),
			fetch              => s_fetch(23,32),
			data_in            => s_data_in(23,32),
			data_out           => s_data_out(23,32),
			out1               => s_out1(23,32),
			out2               => s_out2(23,32),
			lock_lower_row_out => s_locks_lower_out(23,32),
			lock_lower_row_in  => s_locks_lower_in(23,32),
			in1                => s_in1(23,32),
			in2                => s_in2(23,32),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(32)
		);
	s_in1(23,32)            <= s_out1(24,32);
	s_in2(23,32)            <= s_out2(24,33);
	s_locks_lower_in(23,32) <= s_locks_lower_out(24,32);

		normal_cell_23_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,33),
			fetch              => s_fetch(23,33),
			data_in            => s_data_in(23,33),
			data_out           => s_data_out(23,33),
			out1               => s_out1(23,33),
			out2               => s_out2(23,33),
			lock_lower_row_out => s_locks_lower_out(23,33),
			lock_lower_row_in  => s_locks_lower_in(23,33),
			in1                => s_in1(23,33),
			in2                => s_in2(23,33),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(33)
		);
	s_in1(23,33)            <= s_out1(24,33);
	s_in2(23,33)            <= s_out2(24,34);
	s_locks_lower_in(23,33) <= s_locks_lower_out(24,33);

		normal_cell_23_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,34),
			fetch              => s_fetch(23,34),
			data_in            => s_data_in(23,34),
			data_out           => s_data_out(23,34),
			out1               => s_out1(23,34),
			out2               => s_out2(23,34),
			lock_lower_row_out => s_locks_lower_out(23,34),
			lock_lower_row_in  => s_locks_lower_in(23,34),
			in1                => s_in1(23,34),
			in2                => s_in2(23,34),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(34)
		);
	s_in1(23,34)            <= s_out1(24,34);
	s_in2(23,34)            <= s_out2(24,35);
	s_locks_lower_in(23,34) <= s_locks_lower_out(24,34);

		normal_cell_23_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,35),
			fetch              => s_fetch(23,35),
			data_in            => s_data_in(23,35),
			data_out           => s_data_out(23,35),
			out1               => s_out1(23,35),
			out2               => s_out2(23,35),
			lock_lower_row_out => s_locks_lower_out(23,35),
			lock_lower_row_in  => s_locks_lower_in(23,35),
			in1                => s_in1(23,35),
			in2                => s_in2(23,35),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(35)
		);
	s_in1(23,35)            <= s_out1(24,35);
	s_in2(23,35)            <= s_out2(24,36);
	s_locks_lower_in(23,35) <= s_locks_lower_out(24,35);

		normal_cell_23_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,36),
			fetch              => s_fetch(23,36),
			data_in            => s_data_in(23,36),
			data_out           => s_data_out(23,36),
			out1               => s_out1(23,36),
			out2               => s_out2(23,36),
			lock_lower_row_out => s_locks_lower_out(23,36),
			lock_lower_row_in  => s_locks_lower_in(23,36),
			in1                => s_in1(23,36),
			in2                => s_in2(23,36),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(36)
		);
	s_in1(23,36)            <= s_out1(24,36);
	s_in2(23,36)            <= s_out2(24,37);
	s_locks_lower_in(23,36) <= s_locks_lower_out(24,36);

		normal_cell_23_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,37),
			fetch              => s_fetch(23,37),
			data_in            => s_data_in(23,37),
			data_out           => s_data_out(23,37),
			out1               => s_out1(23,37),
			out2               => s_out2(23,37),
			lock_lower_row_out => s_locks_lower_out(23,37),
			lock_lower_row_in  => s_locks_lower_in(23,37),
			in1                => s_in1(23,37),
			in2                => s_in2(23,37),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(37)
		);
	s_in1(23,37)            <= s_out1(24,37);
	s_in2(23,37)            <= s_out2(24,38);
	s_locks_lower_in(23,37) <= s_locks_lower_out(24,37);

		normal_cell_23_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,38),
			fetch              => s_fetch(23,38),
			data_in            => s_data_in(23,38),
			data_out           => s_data_out(23,38),
			out1               => s_out1(23,38),
			out2               => s_out2(23,38),
			lock_lower_row_out => s_locks_lower_out(23,38),
			lock_lower_row_in  => s_locks_lower_in(23,38),
			in1                => s_in1(23,38),
			in2                => s_in2(23,38),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(38)
		);
	s_in1(23,38)            <= s_out1(24,38);
	s_in2(23,38)            <= s_out2(24,39);
	s_locks_lower_in(23,38) <= s_locks_lower_out(24,38);

		normal_cell_23_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,39),
			fetch              => s_fetch(23,39),
			data_in            => s_data_in(23,39),
			data_out           => s_data_out(23,39),
			out1               => s_out1(23,39),
			out2               => s_out2(23,39),
			lock_lower_row_out => s_locks_lower_out(23,39),
			lock_lower_row_in  => s_locks_lower_in(23,39),
			in1                => s_in1(23,39),
			in2                => s_in2(23,39),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(39)
		);
	s_in1(23,39)            <= s_out1(24,39);
	s_in2(23,39)            <= s_out2(24,40);
	s_locks_lower_in(23,39) <= s_locks_lower_out(24,39);

		normal_cell_23_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,40),
			fetch              => s_fetch(23,40),
			data_in            => s_data_in(23,40),
			data_out           => s_data_out(23,40),
			out1               => s_out1(23,40),
			out2               => s_out2(23,40),
			lock_lower_row_out => s_locks_lower_out(23,40),
			lock_lower_row_in  => s_locks_lower_in(23,40),
			in1                => s_in1(23,40),
			in2                => s_in2(23,40),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(40)
		);
	s_in1(23,40)            <= s_out1(24,40);
	s_in2(23,40)            <= s_out2(24,41);
	s_locks_lower_in(23,40) <= s_locks_lower_out(24,40);

		normal_cell_23_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,41),
			fetch              => s_fetch(23,41),
			data_in            => s_data_in(23,41),
			data_out           => s_data_out(23,41),
			out1               => s_out1(23,41),
			out2               => s_out2(23,41),
			lock_lower_row_out => s_locks_lower_out(23,41),
			lock_lower_row_in  => s_locks_lower_in(23,41),
			in1                => s_in1(23,41),
			in2                => s_in2(23,41),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(41)
		);
	s_in1(23,41)            <= s_out1(24,41);
	s_in2(23,41)            <= s_out2(24,42);
	s_locks_lower_in(23,41) <= s_locks_lower_out(24,41);

		normal_cell_23_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,42),
			fetch              => s_fetch(23,42),
			data_in            => s_data_in(23,42),
			data_out           => s_data_out(23,42),
			out1               => s_out1(23,42),
			out2               => s_out2(23,42),
			lock_lower_row_out => s_locks_lower_out(23,42),
			lock_lower_row_in  => s_locks_lower_in(23,42),
			in1                => s_in1(23,42),
			in2                => s_in2(23,42),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(42)
		);
	s_in1(23,42)            <= s_out1(24,42);
	s_in2(23,42)            <= s_out2(24,43);
	s_locks_lower_in(23,42) <= s_locks_lower_out(24,42);

		normal_cell_23_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,43),
			fetch              => s_fetch(23,43),
			data_in            => s_data_in(23,43),
			data_out           => s_data_out(23,43),
			out1               => s_out1(23,43),
			out2               => s_out2(23,43),
			lock_lower_row_out => s_locks_lower_out(23,43),
			lock_lower_row_in  => s_locks_lower_in(23,43),
			in1                => s_in1(23,43),
			in2                => s_in2(23,43),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(43)
		);
	s_in1(23,43)            <= s_out1(24,43);
	s_in2(23,43)            <= s_out2(24,44);
	s_locks_lower_in(23,43) <= s_locks_lower_out(24,43);

		normal_cell_23_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,44),
			fetch              => s_fetch(23,44),
			data_in            => s_data_in(23,44),
			data_out           => s_data_out(23,44),
			out1               => s_out1(23,44),
			out2               => s_out2(23,44),
			lock_lower_row_out => s_locks_lower_out(23,44),
			lock_lower_row_in  => s_locks_lower_in(23,44),
			in1                => s_in1(23,44),
			in2                => s_in2(23,44),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(44)
		);
	s_in1(23,44)            <= s_out1(24,44);
	s_in2(23,44)            <= s_out2(24,45);
	s_locks_lower_in(23,44) <= s_locks_lower_out(24,44);

		normal_cell_23_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,45),
			fetch              => s_fetch(23,45),
			data_in            => s_data_in(23,45),
			data_out           => s_data_out(23,45),
			out1               => s_out1(23,45),
			out2               => s_out2(23,45),
			lock_lower_row_out => s_locks_lower_out(23,45),
			lock_lower_row_in  => s_locks_lower_in(23,45),
			in1                => s_in1(23,45),
			in2                => s_in2(23,45),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(45)
		);
	s_in1(23,45)            <= s_out1(24,45);
	s_in2(23,45)            <= s_out2(24,46);
	s_locks_lower_in(23,45) <= s_locks_lower_out(24,45);

		normal_cell_23_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,46),
			fetch              => s_fetch(23,46),
			data_in            => s_data_in(23,46),
			data_out           => s_data_out(23,46),
			out1               => s_out1(23,46),
			out2               => s_out2(23,46),
			lock_lower_row_out => s_locks_lower_out(23,46),
			lock_lower_row_in  => s_locks_lower_in(23,46),
			in1                => s_in1(23,46),
			in2                => s_in2(23,46),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(46)
		);
	s_in1(23,46)            <= s_out1(24,46);
	s_in2(23,46)            <= s_out2(24,47);
	s_locks_lower_in(23,46) <= s_locks_lower_out(24,46);

		normal_cell_23_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,47),
			fetch              => s_fetch(23,47),
			data_in            => s_data_in(23,47),
			data_out           => s_data_out(23,47),
			out1               => s_out1(23,47),
			out2               => s_out2(23,47),
			lock_lower_row_out => s_locks_lower_out(23,47),
			lock_lower_row_in  => s_locks_lower_in(23,47),
			in1                => s_in1(23,47),
			in2                => s_in2(23,47),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(47)
		);
	s_in1(23,47)            <= s_out1(24,47);
	s_in2(23,47)            <= s_out2(24,48);
	s_locks_lower_in(23,47) <= s_locks_lower_out(24,47);

		normal_cell_23_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,48),
			fetch              => s_fetch(23,48),
			data_in            => s_data_in(23,48),
			data_out           => s_data_out(23,48),
			out1               => s_out1(23,48),
			out2               => s_out2(23,48),
			lock_lower_row_out => s_locks_lower_out(23,48),
			lock_lower_row_in  => s_locks_lower_in(23,48),
			in1                => s_in1(23,48),
			in2                => s_in2(23,48),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(48)
		);
	s_in1(23,48)            <= s_out1(24,48);
	s_in2(23,48)            <= s_out2(24,49);
	s_locks_lower_in(23,48) <= s_locks_lower_out(24,48);

		normal_cell_23_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,49),
			fetch              => s_fetch(23,49),
			data_in            => s_data_in(23,49),
			data_out           => s_data_out(23,49),
			out1               => s_out1(23,49),
			out2               => s_out2(23,49),
			lock_lower_row_out => s_locks_lower_out(23,49),
			lock_lower_row_in  => s_locks_lower_in(23,49),
			in1                => s_in1(23,49),
			in2                => s_in2(23,49),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(49)
		);
	s_in1(23,49)            <= s_out1(24,49);
	s_in2(23,49)            <= s_out2(24,50);
	s_locks_lower_in(23,49) <= s_locks_lower_out(24,49);

		normal_cell_23_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,50),
			fetch              => s_fetch(23,50),
			data_in            => s_data_in(23,50),
			data_out           => s_data_out(23,50),
			out1               => s_out1(23,50),
			out2               => s_out2(23,50),
			lock_lower_row_out => s_locks_lower_out(23,50),
			lock_lower_row_in  => s_locks_lower_in(23,50),
			in1                => s_in1(23,50),
			in2                => s_in2(23,50),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(50)
		);
	s_in1(23,50)            <= s_out1(24,50);
	s_in2(23,50)            <= s_out2(24,51);
	s_locks_lower_in(23,50) <= s_locks_lower_out(24,50);

		normal_cell_23_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,51),
			fetch              => s_fetch(23,51),
			data_in            => s_data_in(23,51),
			data_out           => s_data_out(23,51),
			out1               => s_out1(23,51),
			out2               => s_out2(23,51),
			lock_lower_row_out => s_locks_lower_out(23,51),
			lock_lower_row_in  => s_locks_lower_in(23,51),
			in1                => s_in1(23,51),
			in2                => s_in2(23,51),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(51)
		);
	s_in1(23,51)            <= s_out1(24,51);
	s_in2(23,51)            <= s_out2(24,52);
	s_locks_lower_in(23,51) <= s_locks_lower_out(24,51);

		normal_cell_23_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,52),
			fetch              => s_fetch(23,52),
			data_in            => s_data_in(23,52),
			data_out           => s_data_out(23,52),
			out1               => s_out1(23,52),
			out2               => s_out2(23,52),
			lock_lower_row_out => s_locks_lower_out(23,52),
			lock_lower_row_in  => s_locks_lower_in(23,52),
			in1                => s_in1(23,52),
			in2                => s_in2(23,52),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(52)
		);
	s_in1(23,52)            <= s_out1(24,52);
	s_in2(23,52)            <= s_out2(24,53);
	s_locks_lower_in(23,52) <= s_locks_lower_out(24,52);

		normal_cell_23_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,53),
			fetch              => s_fetch(23,53),
			data_in            => s_data_in(23,53),
			data_out           => s_data_out(23,53),
			out1               => s_out1(23,53),
			out2               => s_out2(23,53),
			lock_lower_row_out => s_locks_lower_out(23,53),
			lock_lower_row_in  => s_locks_lower_in(23,53),
			in1                => s_in1(23,53),
			in2                => s_in2(23,53),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(53)
		);
	s_in1(23,53)            <= s_out1(24,53);
	s_in2(23,53)            <= s_out2(24,54);
	s_locks_lower_in(23,53) <= s_locks_lower_out(24,53);

		normal_cell_23_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,54),
			fetch              => s_fetch(23,54),
			data_in            => s_data_in(23,54),
			data_out           => s_data_out(23,54),
			out1               => s_out1(23,54),
			out2               => s_out2(23,54),
			lock_lower_row_out => s_locks_lower_out(23,54),
			lock_lower_row_in  => s_locks_lower_in(23,54),
			in1                => s_in1(23,54),
			in2                => s_in2(23,54),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(54)
		);
	s_in1(23,54)            <= s_out1(24,54);
	s_in2(23,54)            <= s_out2(24,55);
	s_locks_lower_in(23,54) <= s_locks_lower_out(24,54);

		normal_cell_23_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,55),
			fetch              => s_fetch(23,55),
			data_in            => s_data_in(23,55),
			data_out           => s_data_out(23,55),
			out1               => s_out1(23,55),
			out2               => s_out2(23,55),
			lock_lower_row_out => s_locks_lower_out(23,55),
			lock_lower_row_in  => s_locks_lower_in(23,55),
			in1                => s_in1(23,55),
			in2                => s_in2(23,55),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(55)
		);
	s_in1(23,55)            <= s_out1(24,55);
	s_in2(23,55)            <= s_out2(24,56);
	s_locks_lower_in(23,55) <= s_locks_lower_out(24,55);

		normal_cell_23_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,56),
			fetch              => s_fetch(23,56),
			data_in            => s_data_in(23,56),
			data_out           => s_data_out(23,56),
			out1               => s_out1(23,56),
			out2               => s_out2(23,56),
			lock_lower_row_out => s_locks_lower_out(23,56),
			lock_lower_row_in  => s_locks_lower_in(23,56),
			in1                => s_in1(23,56),
			in2                => s_in2(23,56),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(56)
		);
	s_in1(23,56)            <= s_out1(24,56);
	s_in2(23,56)            <= s_out2(24,57);
	s_locks_lower_in(23,56) <= s_locks_lower_out(24,56);

		normal_cell_23_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,57),
			fetch              => s_fetch(23,57),
			data_in            => s_data_in(23,57),
			data_out           => s_data_out(23,57),
			out1               => s_out1(23,57),
			out2               => s_out2(23,57),
			lock_lower_row_out => s_locks_lower_out(23,57),
			lock_lower_row_in  => s_locks_lower_in(23,57),
			in1                => s_in1(23,57),
			in2                => s_in2(23,57),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(57)
		);
	s_in1(23,57)            <= s_out1(24,57);
	s_in2(23,57)            <= s_out2(24,58);
	s_locks_lower_in(23,57) <= s_locks_lower_out(24,57);

		normal_cell_23_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,58),
			fetch              => s_fetch(23,58),
			data_in            => s_data_in(23,58),
			data_out           => s_data_out(23,58),
			out1               => s_out1(23,58),
			out2               => s_out2(23,58),
			lock_lower_row_out => s_locks_lower_out(23,58),
			lock_lower_row_in  => s_locks_lower_in(23,58),
			in1                => s_in1(23,58),
			in2                => s_in2(23,58),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(58)
		);
	s_in1(23,58)            <= s_out1(24,58);
	s_in2(23,58)            <= s_out2(24,59);
	s_locks_lower_in(23,58) <= s_locks_lower_out(24,58);

		normal_cell_23_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,59),
			fetch              => s_fetch(23,59),
			data_in            => s_data_in(23,59),
			data_out           => s_data_out(23,59),
			out1               => s_out1(23,59),
			out2               => s_out2(23,59),
			lock_lower_row_out => s_locks_lower_out(23,59),
			lock_lower_row_in  => s_locks_lower_in(23,59),
			in1                => s_in1(23,59),
			in2                => s_in2(23,59),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(59)
		);
	s_in1(23,59)            <= s_out1(24,59);
	s_in2(23,59)            <= s_out2(24,60);
	s_locks_lower_in(23,59) <= s_locks_lower_out(24,59);

		last_col_cell_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(23,60),
			fetch              => s_fetch(23,60),
			data_in            => s_data_in(23,60),
			data_out           => s_data_out(23,60),
			out1               => s_out1(23,60),
			out2               => s_out2(23,60),
			lock_lower_row_out => s_locks_lower_out(23,60),
			lock_lower_row_in  => s_locks_lower_in(23,60),
			in1                => s_in1(23,60),
			in2                => (others => '0'),
			lock_row           => s_locks(23),
			piv_found          => s_piv_found,
			row_data           => s_row_data(23),
			col_data           => s_col_data(60)
		);
	s_in1(23,60)            <= s_out1(24,60);
	s_locks_lower_in(23,60) <= s_locks_lower_out(24,60);

		normal_cell_24_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,1),
			fetch              => s_fetch(24,1),
			data_in            => s_data_in(24,1),
			data_out           => s_data_out(24,1),
			out1               => s_out1(24,1),
			out2               => s_out2(24,1),
			lock_lower_row_out => s_locks_lower_out(24,1),
			lock_lower_row_in  => s_locks_lower_in(24,1),
			in1                => s_in1(24,1),
			in2                => s_in2(24,1),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(1)
		);
	s_in1(24,1)            <= s_out1(25,1);
	s_in2(24,1)            <= s_out2(25,2);
	s_locks_lower_in(24,1) <= s_locks_lower_out(25,1);

		normal_cell_24_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,2),
			fetch              => s_fetch(24,2),
			data_in            => s_data_in(24,2),
			data_out           => s_data_out(24,2),
			out1               => s_out1(24,2),
			out2               => s_out2(24,2),
			lock_lower_row_out => s_locks_lower_out(24,2),
			lock_lower_row_in  => s_locks_lower_in(24,2),
			in1                => s_in1(24,2),
			in2                => s_in2(24,2),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(2)
		);
	s_in1(24,2)            <= s_out1(25,2);
	s_in2(24,2)            <= s_out2(25,3);
	s_locks_lower_in(24,2) <= s_locks_lower_out(25,2);

		normal_cell_24_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,3),
			fetch              => s_fetch(24,3),
			data_in            => s_data_in(24,3),
			data_out           => s_data_out(24,3),
			out1               => s_out1(24,3),
			out2               => s_out2(24,3),
			lock_lower_row_out => s_locks_lower_out(24,3),
			lock_lower_row_in  => s_locks_lower_in(24,3),
			in1                => s_in1(24,3),
			in2                => s_in2(24,3),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(3)
		);
	s_in1(24,3)            <= s_out1(25,3);
	s_in2(24,3)            <= s_out2(25,4);
	s_locks_lower_in(24,3) <= s_locks_lower_out(25,3);

		normal_cell_24_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,4),
			fetch              => s_fetch(24,4),
			data_in            => s_data_in(24,4),
			data_out           => s_data_out(24,4),
			out1               => s_out1(24,4),
			out2               => s_out2(24,4),
			lock_lower_row_out => s_locks_lower_out(24,4),
			lock_lower_row_in  => s_locks_lower_in(24,4),
			in1                => s_in1(24,4),
			in2                => s_in2(24,4),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(4)
		);
	s_in1(24,4)            <= s_out1(25,4);
	s_in2(24,4)            <= s_out2(25,5);
	s_locks_lower_in(24,4) <= s_locks_lower_out(25,4);

		normal_cell_24_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,5),
			fetch              => s_fetch(24,5),
			data_in            => s_data_in(24,5),
			data_out           => s_data_out(24,5),
			out1               => s_out1(24,5),
			out2               => s_out2(24,5),
			lock_lower_row_out => s_locks_lower_out(24,5),
			lock_lower_row_in  => s_locks_lower_in(24,5),
			in1                => s_in1(24,5),
			in2                => s_in2(24,5),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(5)
		);
	s_in1(24,5)            <= s_out1(25,5);
	s_in2(24,5)            <= s_out2(25,6);
	s_locks_lower_in(24,5) <= s_locks_lower_out(25,5);

		normal_cell_24_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,6),
			fetch              => s_fetch(24,6),
			data_in            => s_data_in(24,6),
			data_out           => s_data_out(24,6),
			out1               => s_out1(24,6),
			out2               => s_out2(24,6),
			lock_lower_row_out => s_locks_lower_out(24,6),
			lock_lower_row_in  => s_locks_lower_in(24,6),
			in1                => s_in1(24,6),
			in2                => s_in2(24,6),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(6)
		);
	s_in1(24,6)            <= s_out1(25,6);
	s_in2(24,6)            <= s_out2(25,7);
	s_locks_lower_in(24,6) <= s_locks_lower_out(25,6);

		normal_cell_24_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,7),
			fetch              => s_fetch(24,7),
			data_in            => s_data_in(24,7),
			data_out           => s_data_out(24,7),
			out1               => s_out1(24,7),
			out2               => s_out2(24,7),
			lock_lower_row_out => s_locks_lower_out(24,7),
			lock_lower_row_in  => s_locks_lower_in(24,7),
			in1                => s_in1(24,7),
			in2                => s_in2(24,7),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(7)
		);
	s_in1(24,7)            <= s_out1(25,7);
	s_in2(24,7)            <= s_out2(25,8);
	s_locks_lower_in(24,7) <= s_locks_lower_out(25,7);

		normal_cell_24_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,8),
			fetch              => s_fetch(24,8),
			data_in            => s_data_in(24,8),
			data_out           => s_data_out(24,8),
			out1               => s_out1(24,8),
			out2               => s_out2(24,8),
			lock_lower_row_out => s_locks_lower_out(24,8),
			lock_lower_row_in  => s_locks_lower_in(24,8),
			in1                => s_in1(24,8),
			in2                => s_in2(24,8),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(8)
		);
	s_in1(24,8)            <= s_out1(25,8);
	s_in2(24,8)            <= s_out2(25,9);
	s_locks_lower_in(24,8) <= s_locks_lower_out(25,8);

		normal_cell_24_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,9),
			fetch              => s_fetch(24,9),
			data_in            => s_data_in(24,9),
			data_out           => s_data_out(24,9),
			out1               => s_out1(24,9),
			out2               => s_out2(24,9),
			lock_lower_row_out => s_locks_lower_out(24,9),
			lock_lower_row_in  => s_locks_lower_in(24,9),
			in1                => s_in1(24,9),
			in2                => s_in2(24,9),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(9)
		);
	s_in1(24,9)            <= s_out1(25,9);
	s_in2(24,9)            <= s_out2(25,10);
	s_locks_lower_in(24,9) <= s_locks_lower_out(25,9);

		normal_cell_24_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,10),
			fetch              => s_fetch(24,10),
			data_in            => s_data_in(24,10),
			data_out           => s_data_out(24,10),
			out1               => s_out1(24,10),
			out2               => s_out2(24,10),
			lock_lower_row_out => s_locks_lower_out(24,10),
			lock_lower_row_in  => s_locks_lower_in(24,10),
			in1                => s_in1(24,10),
			in2                => s_in2(24,10),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(10)
		);
	s_in1(24,10)            <= s_out1(25,10);
	s_in2(24,10)            <= s_out2(25,11);
	s_locks_lower_in(24,10) <= s_locks_lower_out(25,10);

		normal_cell_24_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,11),
			fetch              => s_fetch(24,11),
			data_in            => s_data_in(24,11),
			data_out           => s_data_out(24,11),
			out1               => s_out1(24,11),
			out2               => s_out2(24,11),
			lock_lower_row_out => s_locks_lower_out(24,11),
			lock_lower_row_in  => s_locks_lower_in(24,11),
			in1                => s_in1(24,11),
			in2                => s_in2(24,11),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(11)
		);
	s_in1(24,11)            <= s_out1(25,11);
	s_in2(24,11)            <= s_out2(25,12);
	s_locks_lower_in(24,11) <= s_locks_lower_out(25,11);

		normal_cell_24_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,12),
			fetch              => s_fetch(24,12),
			data_in            => s_data_in(24,12),
			data_out           => s_data_out(24,12),
			out1               => s_out1(24,12),
			out2               => s_out2(24,12),
			lock_lower_row_out => s_locks_lower_out(24,12),
			lock_lower_row_in  => s_locks_lower_in(24,12),
			in1                => s_in1(24,12),
			in2                => s_in2(24,12),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(12)
		);
	s_in1(24,12)            <= s_out1(25,12);
	s_in2(24,12)            <= s_out2(25,13);
	s_locks_lower_in(24,12) <= s_locks_lower_out(25,12);

		normal_cell_24_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,13),
			fetch              => s_fetch(24,13),
			data_in            => s_data_in(24,13),
			data_out           => s_data_out(24,13),
			out1               => s_out1(24,13),
			out2               => s_out2(24,13),
			lock_lower_row_out => s_locks_lower_out(24,13),
			lock_lower_row_in  => s_locks_lower_in(24,13),
			in1                => s_in1(24,13),
			in2                => s_in2(24,13),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(13)
		);
	s_in1(24,13)            <= s_out1(25,13);
	s_in2(24,13)            <= s_out2(25,14);
	s_locks_lower_in(24,13) <= s_locks_lower_out(25,13);

		normal_cell_24_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,14),
			fetch              => s_fetch(24,14),
			data_in            => s_data_in(24,14),
			data_out           => s_data_out(24,14),
			out1               => s_out1(24,14),
			out2               => s_out2(24,14),
			lock_lower_row_out => s_locks_lower_out(24,14),
			lock_lower_row_in  => s_locks_lower_in(24,14),
			in1                => s_in1(24,14),
			in2                => s_in2(24,14),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(14)
		);
	s_in1(24,14)            <= s_out1(25,14);
	s_in2(24,14)            <= s_out2(25,15);
	s_locks_lower_in(24,14) <= s_locks_lower_out(25,14);

		normal_cell_24_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,15),
			fetch              => s_fetch(24,15),
			data_in            => s_data_in(24,15),
			data_out           => s_data_out(24,15),
			out1               => s_out1(24,15),
			out2               => s_out2(24,15),
			lock_lower_row_out => s_locks_lower_out(24,15),
			lock_lower_row_in  => s_locks_lower_in(24,15),
			in1                => s_in1(24,15),
			in2                => s_in2(24,15),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(15)
		);
	s_in1(24,15)            <= s_out1(25,15);
	s_in2(24,15)            <= s_out2(25,16);
	s_locks_lower_in(24,15) <= s_locks_lower_out(25,15);

		normal_cell_24_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,16),
			fetch              => s_fetch(24,16),
			data_in            => s_data_in(24,16),
			data_out           => s_data_out(24,16),
			out1               => s_out1(24,16),
			out2               => s_out2(24,16),
			lock_lower_row_out => s_locks_lower_out(24,16),
			lock_lower_row_in  => s_locks_lower_in(24,16),
			in1                => s_in1(24,16),
			in2                => s_in2(24,16),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(16)
		);
	s_in1(24,16)            <= s_out1(25,16);
	s_in2(24,16)            <= s_out2(25,17);
	s_locks_lower_in(24,16) <= s_locks_lower_out(25,16);

		normal_cell_24_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,17),
			fetch              => s_fetch(24,17),
			data_in            => s_data_in(24,17),
			data_out           => s_data_out(24,17),
			out1               => s_out1(24,17),
			out2               => s_out2(24,17),
			lock_lower_row_out => s_locks_lower_out(24,17),
			lock_lower_row_in  => s_locks_lower_in(24,17),
			in1                => s_in1(24,17),
			in2                => s_in2(24,17),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(17)
		);
	s_in1(24,17)            <= s_out1(25,17);
	s_in2(24,17)            <= s_out2(25,18);
	s_locks_lower_in(24,17) <= s_locks_lower_out(25,17);

		normal_cell_24_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,18),
			fetch              => s_fetch(24,18),
			data_in            => s_data_in(24,18),
			data_out           => s_data_out(24,18),
			out1               => s_out1(24,18),
			out2               => s_out2(24,18),
			lock_lower_row_out => s_locks_lower_out(24,18),
			lock_lower_row_in  => s_locks_lower_in(24,18),
			in1                => s_in1(24,18),
			in2                => s_in2(24,18),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(18)
		);
	s_in1(24,18)            <= s_out1(25,18);
	s_in2(24,18)            <= s_out2(25,19);
	s_locks_lower_in(24,18) <= s_locks_lower_out(25,18);

		normal_cell_24_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,19),
			fetch              => s_fetch(24,19),
			data_in            => s_data_in(24,19),
			data_out           => s_data_out(24,19),
			out1               => s_out1(24,19),
			out2               => s_out2(24,19),
			lock_lower_row_out => s_locks_lower_out(24,19),
			lock_lower_row_in  => s_locks_lower_in(24,19),
			in1                => s_in1(24,19),
			in2                => s_in2(24,19),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(19)
		);
	s_in1(24,19)            <= s_out1(25,19);
	s_in2(24,19)            <= s_out2(25,20);
	s_locks_lower_in(24,19) <= s_locks_lower_out(25,19);

		normal_cell_24_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,20),
			fetch              => s_fetch(24,20),
			data_in            => s_data_in(24,20),
			data_out           => s_data_out(24,20),
			out1               => s_out1(24,20),
			out2               => s_out2(24,20),
			lock_lower_row_out => s_locks_lower_out(24,20),
			lock_lower_row_in  => s_locks_lower_in(24,20),
			in1                => s_in1(24,20),
			in2                => s_in2(24,20),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(20)
		);
	s_in1(24,20)            <= s_out1(25,20);
	s_in2(24,20)            <= s_out2(25,21);
	s_locks_lower_in(24,20) <= s_locks_lower_out(25,20);

		normal_cell_24_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,21),
			fetch              => s_fetch(24,21),
			data_in            => s_data_in(24,21),
			data_out           => s_data_out(24,21),
			out1               => s_out1(24,21),
			out2               => s_out2(24,21),
			lock_lower_row_out => s_locks_lower_out(24,21),
			lock_lower_row_in  => s_locks_lower_in(24,21),
			in1                => s_in1(24,21),
			in2                => s_in2(24,21),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(21)
		);
	s_in1(24,21)            <= s_out1(25,21);
	s_in2(24,21)            <= s_out2(25,22);
	s_locks_lower_in(24,21) <= s_locks_lower_out(25,21);

		normal_cell_24_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,22),
			fetch              => s_fetch(24,22),
			data_in            => s_data_in(24,22),
			data_out           => s_data_out(24,22),
			out1               => s_out1(24,22),
			out2               => s_out2(24,22),
			lock_lower_row_out => s_locks_lower_out(24,22),
			lock_lower_row_in  => s_locks_lower_in(24,22),
			in1                => s_in1(24,22),
			in2                => s_in2(24,22),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(22)
		);
	s_in1(24,22)            <= s_out1(25,22);
	s_in2(24,22)            <= s_out2(25,23);
	s_locks_lower_in(24,22) <= s_locks_lower_out(25,22);

		normal_cell_24_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,23),
			fetch              => s_fetch(24,23),
			data_in            => s_data_in(24,23),
			data_out           => s_data_out(24,23),
			out1               => s_out1(24,23),
			out2               => s_out2(24,23),
			lock_lower_row_out => s_locks_lower_out(24,23),
			lock_lower_row_in  => s_locks_lower_in(24,23),
			in1                => s_in1(24,23),
			in2                => s_in2(24,23),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(23)
		);
	s_in1(24,23)            <= s_out1(25,23);
	s_in2(24,23)            <= s_out2(25,24);
	s_locks_lower_in(24,23) <= s_locks_lower_out(25,23);

		normal_cell_24_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,24),
			fetch              => s_fetch(24,24),
			data_in            => s_data_in(24,24),
			data_out           => s_data_out(24,24),
			out1               => s_out1(24,24),
			out2               => s_out2(24,24),
			lock_lower_row_out => s_locks_lower_out(24,24),
			lock_lower_row_in  => s_locks_lower_in(24,24),
			in1                => s_in1(24,24),
			in2                => s_in2(24,24),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(24)
		);
	s_in1(24,24)            <= s_out1(25,24);
	s_in2(24,24)            <= s_out2(25,25);
	s_locks_lower_in(24,24) <= s_locks_lower_out(25,24);

		normal_cell_24_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,25),
			fetch              => s_fetch(24,25),
			data_in            => s_data_in(24,25),
			data_out           => s_data_out(24,25),
			out1               => s_out1(24,25),
			out2               => s_out2(24,25),
			lock_lower_row_out => s_locks_lower_out(24,25),
			lock_lower_row_in  => s_locks_lower_in(24,25),
			in1                => s_in1(24,25),
			in2                => s_in2(24,25),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(25)
		);
	s_in1(24,25)            <= s_out1(25,25);
	s_in2(24,25)            <= s_out2(25,26);
	s_locks_lower_in(24,25) <= s_locks_lower_out(25,25);

		normal_cell_24_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,26),
			fetch              => s_fetch(24,26),
			data_in            => s_data_in(24,26),
			data_out           => s_data_out(24,26),
			out1               => s_out1(24,26),
			out2               => s_out2(24,26),
			lock_lower_row_out => s_locks_lower_out(24,26),
			lock_lower_row_in  => s_locks_lower_in(24,26),
			in1                => s_in1(24,26),
			in2                => s_in2(24,26),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(26)
		);
	s_in1(24,26)            <= s_out1(25,26);
	s_in2(24,26)            <= s_out2(25,27);
	s_locks_lower_in(24,26) <= s_locks_lower_out(25,26);

		normal_cell_24_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,27),
			fetch              => s_fetch(24,27),
			data_in            => s_data_in(24,27),
			data_out           => s_data_out(24,27),
			out1               => s_out1(24,27),
			out2               => s_out2(24,27),
			lock_lower_row_out => s_locks_lower_out(24,27),
			lock_lower_row_in  => s_locks_lower_in(24,27),
			in1                => s_in1(24,27),
			in2                => s_in2(24,27),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(27)
		);
	s_in1(24,27)            <= s_out1(25,27);
	s_in2(24,27)            <= s_out2(25,28);
	s_locks_lower_in(24,27) <= s_locks_lower_out(25,27);

		normal_cell_24_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,28),
			fetch              => s_fetch(24,28),
			data_in            => s_data_in(24,28),
			data_out           => s_data_out(24,28),
			out1               => s_out1(24,28),
			out2               => s_out2(24,28),
			lock_lower_row_out => s_locks_lower_out(24,28),
			lock_lower_row_in  => s_locks_lower_in(24,28),
			in1                => s_in1(24,28),
			in2                => s_in2(24,28),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(28)
		);
	s_in1(24,28)            <= s_out1(25,28);
	s_in2(24,28)            <= s_out2(25,29);
	s_locks_lower_in(24,28) <= s_locks_lower_out(25,28);

		normal_cell_24_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,29),
			fetch              => s_fetch(24,29),
			data_in            => s_data_in(24,29),
			data_out           => s_data_out(24,29),
			out1               => s_out1(24,29),
			out2               => s_out2(24,29),
			lock_lower_row_out => s_locks_lower_out(24,29),
			lock_lower_row_in  => s_locks_lower_in(24,29),
			in1                => s_in1(24,29),
			in2                => s_in2(24,29),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(29)
		);
	s_in1(24,29)            <= s_out1(25,29);
	s_in2(24,29)            <= s_out2(25,30);
	s_locks_lower_in(24,29) <= s_locks_lower_out(25,29);

		normal_cell_24_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,30),
			fetch              => s_fetch(24,30),
			data_in            => s_data_in(24,30),
			data_out           => s_data_out(24,30),
			out1               => s_out1(24,30),
			out2               => s_out2(24,30),
			lock_lower_row_out => s_locks_lower_out(24,30),
			lock_lower_row_in  => s_locks_lower_in(24,30),
			in1                => s_in1(24,30),
			in2                => s_in2(24,30),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(30)
		);
	s_in1(24,30)            <= s_out1(25,30);
	s_in2(24,30)            <= s_out2(25,31);
	s_locks_lower_in(24,30) <= s_locks_lower_out(25,30);

		normal_cell_24_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,31),
			fetch              => s_fetch(24,31),
			data_in            => s_data_in(24,31),
			data_out           => s_data_out(24,31),
			out1               => s_out1(24,31),
			out2               => s_out2(24,31),
			lock_lower_row_out => s_locks_lower_out(24,31),
			lock_lower_row_in  => s_locks_lower_in(24,31),
			in1                => s_in1(24,31),
			in2                => s_in2(24,31),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(31)
		);
	s_in1(24,31)            <= s_out1(25,31);
	s_in2(24,31)            <= s_out2(25,32);
	s_locks_lower_in(24,31) <= s_locks_lower_out(25,31);

		normal_cell_24_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,32),
			fetch              => s_fetch(24,32),
			data_in            => s_data_in(24,32),
			data_out           => s_data_out(24,32),
			out1               => s_out1(24,32),
			out2               => s_out2(24,32),
			lock_lower_row_out => s_locks_lower_out(24,32),
			lock_lower_row_in  => s_locks_lower_in(24,32),
			in1                => s_in1(24,32),
			in2                => s_in2(24,32),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(32)
		);
	s_in1(24,32)            <= s_out1(25,32);
	s_in2(24,32)            <= s_out2(25,33);
	s_locks_lower_in(24,32) <= s_locks_lower_out(25,32);

		normal_cell_24_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,33),
			fetch              => s_fetch(24,33),
			data_in            => s_data_in(24,33),
			data_out           => s_data_out(24,33),
			out1               => s_out1(24,33),
			out2               => s_out2(24,33),
			lock_lower_row_out => s_locks_lower_out(24,33),
			lock_lower_row_in  => s_locks_lower_in(24,33),
			in1                => s_in1(24,33),
			in2                => s_in2(24,33),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(33)
		);
	s_in1(24,33)            <= s_out1(25,33);
	s_in2(24,33)            <= s_out2(25,34);
	s_locks_lower_in(24,33) <= s_locks_lower_out(25,33);

		normal_cell_24_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,34),
			fetch              => s_fetch(24,34),
			data_in            => s_data_in(24,34),
			data_out           => s_data_out(24,34),
			out1               => s_out1(24,34),
			out2               => s_out2(24,34),
			lock_lower_row_out => s_locks_lower_out(24,34),
			lock_lower_row_in  => s_locks_lower_in(24,34),
			in1                => s_in1(24,34),
			in2                => s_in2(24,34),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(34)
		);
	s_in1(24,34)            <= s_out1(25,34);
	s_in2(24,34)            <= s_out2(25,35);
	s_locks_lower_in(24,34) <= s_locks_lower_out(25,34);

		normal_cell_24_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,35),
			fetch              => s_fetch(24,35),
			data_in            => s_data_in(24,35),
			data_out           => s_data_out(24,35),
			out1               => s_out1(24,35),
			out2               => s_out2(24,35),
			lock_lower_row_out => s_locks_lower_out(24,35),
			lock_lower_row_in  => s_locks_lower_in(24,35),
			in1                => s_in1(24,35),
			in2                => s_in2(24,35),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(35)
		);
	s_in1(24,35)            <= s_out1(25,35);
	s_in2(24,35)            <= s_out2(25,36);
	s_locks_lower_in(24,35) <= s_locks_lower_out(25,35);

		normal_cell_24_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,36),
			fetch              => s_fetch(24,36),
			data_in            => s_data_in(24,36),
			data_out           => s_data_out(24,36),
			out1               => s_out1(24,36),
			out2               => s_out2(24,36),
			lock_lower_row_out => s_locks_lower_out(24,36),
			lock_lower_row_in  => s_locks_lower_in(24,36),
			in1                => s_in1(24,36),
			in2                => s_in2(24,36),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(36)
		);
	s_in1(24,36)            <= s_out1(25,36);
	s_in2(24,36)            <= s_out2(25,37);
	s_locks_lower_in(24,36) <= s_locks_lower_out(25,36);

		normal_cell_24_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,37),
			fetch              => s_fetch(24,37),
			data_in            => s_data_in(24,37),
			data_out           => s_data_out(24,37),
			out1               => s_out1(24,37),
			out2               => s_out2(24,37),
			lock_lower_row_out => s_locks_lower_out(24,37),
			lock_lower_row_in  => s_locks_lower_in(24,37),
			in1                => s_in1(24,37),
			in2                => s_in2(24,37),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(37)
		);
	s_in1(24,37)            <= s_out1(25,37);
	s_in2(24,37)            <= s_out2(25,38);
	s_locks_lower_in(24,37) <= s_locks_lower_out(25,37);

		normal_cell_24_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,38),
			fetch              => s_fetch(24,38),
			data_in            => s_data_in(24,38),
			data_out           => s_data_out(24,38),
			out1               => s_out1(24,38),
			out2               => s_out2(24,38),
			lock_lower_row_out => s_locks_lower_out(24,38),
			lock_lower_row_in  => s_locks_lower_in(24,38),
			in1                => s_in1(24,38),
			in2                => s_in2(24,38),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(38)
		);
	s_in1(24,38)            <= s_out1(25,38);
	s_in2(24,38)            <= s_out2(25,39);
	s_locks_lower_in(24,38) <= s_locks_lower_out(25,38);

		normal_cell_24_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,39),
			fetch              => s_fetch(24,39),
			data_in            => s_data_in(24,39),
			data_out           => s_data_out(24,39),
			out1               => s_out1(24,39),
			out2               => s_out2(24,39),
			lock_lower_row_out => s_locks_lower_out(24,39),
			lock_lower_row_in  => s_locks_lower_in(24,39),
			in1                => s_in1(24,39),
			in2                => s_in2(24,39),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(39)
		);
	s_in1(24,39)            <= s_out1(25,39);
	s_in2(24,39)            <= s_out2(25,40);
	s_locks_lower_in(24,39) <= s_locks_lower_out(25,39);

		normal_cell_24_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,40),
			fetch              => s_fetch(24,40),
			data_in            => s_data_in(24,40),
			data_out           => s_data_out(24,40),
			out1               => s_out1(24,40),
			out2               => s_out2(24,40),
			lock_lower_row_out => s_locks_lower_out(24,40),
			lock_lower_row_in  => s_locks_lower_in(24,40),
			in1                => s_in1(24,40),
			in2                => s_in2(24,40),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(40)
		);
	s_in1(24,40)            <= s_out1(25,40);
	s_in2(24,40)            <= s_out2(25,41);
	s_locks_lower_in(24,40) <= s_locks_lower_out(25,40);

		normal_cell_24_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,41),
			fetch              => s_fetch(24,41),
			data_in            => s_data_in(24,41),
			data_out           => s_data_out(24,41),
			out1               => s_out1(24,41),
			out2               => s_out2(24,41),
			lock_lower_row_out => s_locks_lower_out(24,41),
			lock_lower_row_in  => s_locks_lower_in(24,41),
			in1                => s_in1(24,41),
			in2                => s_in2(24,41),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(41)
		);
	s_in1(24,41)            <= s_out1(25,41);
	s_in2(24,41)            <= s_out2(25,42);
	s_locks_lower_in(24,41) <= s_locks_lower_out(25,41);

		normal_cell_24_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,42),
			fetch              => s_fetch(24,42),
			data_in            => s_data_in(24,42),
			data_out           => s_data_out(24,42),
			out1               => s_out1(24,42),
			out2               => s_out2(24,42),
			lock_lower_row_out => s_locks_lower_out(24,42),
			lock_lower_row_in  => s_locks_lower_in(24,42),
			in1                => s_in1(24,42),
			in2                => s_in2(24,42),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(42)
		);
	s_in1(24,42)            <= s_out1(25,42);
	s_in2(24,42)            <= s_out2(25,43);
	s_locks_lower_in(24,42) <= s_locks_lower_out(25,42);

		normal_cell_24_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,43),
			fetch              => s_fetch(24,43),
			data_in            => s_data_in(24,43),
			data_out           => s_data_out(24,43),
			out1               => s_out1(24,43),
			out2               => s_out2(24,43),
			lock_lower_row_out => s_locks_lower_out(24,43),
			lock_lower_row_in  => s_locks_lower_in(24,43),
			in1                => s_in1(24,43),
			in2                => s_in2(24,43),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(43)
		);
	s_in1(24,43)            <= s_out1(25,43);
	s_in2(24,43)            <= s_out2(25,44);
	s_locks_lower_in(24,43) <= s_locks_lower_out(25,43);

		normal_cell_24_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,44),
			fetch              => s_fetch(24,44),
			data_in            => s_data_in(24,44),
			data_out           => s_data_out(24,44),
			out1               => s_out1(24,44),
			out2               => s_out2(24,44),
			lock_lower_row_out => s_locks_lower_out(24,44),
			lock_lower_row_in  => s_locks_lower_in(24,44),
			in1                => s_in1(24,44),
			in2                => s_in2(24,44),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(44)
		);
	s_in1(24,44)            <= s_out1(25,44);
	s_in2(24,44)            <= s_out2(25,45);
	s_locks_lower_in(24,44) <= s_locks_lower_out(25,44);

		normal_cell_24_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,45),
			fetch              => s_fetch(24,45),
			data_in            => s_data_in(24,45),
			data_out           => s_data_out(24,45),
			out1               => s_out1(24,45),
			out2               => s_out2(24,45),
			lock_lower_row_out => s_locks_lower_out(24,45),
			lock_lower_row_in  => s_locks_lower_in(24,45),
			in1                => s_in1(24,45),
			in2                => s_in2(24,45),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(45)
		);
	s_in1(24,45)            <= s_out1(25,45);
	s_in2(24,45)            <= s_out2(25,46);
	s_locks_lower_in(24,45) <= s_locks_lower_out(25,45);

		normal_cell_24_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,46),
			fetch              => s_fetch(24,46),
			data_in            => s_data_in(24,46),
			data_out           => s_data_out(24,46),
			out1               => s_out1(24,46),
			out2               => s_out2(24,46),
			lock_lower_row_out => s_locks_lower_out(24,46),
			lock_lower_row_in  => s_locks_lower_in(24,46),
			in1                => s_in1(24,46),
			in2                => s_in2(24,46),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(46)
		);
	s_in1(24,46)            <= s_out1(25,46);
	s_in2(24,46)            <= s_out2(25,47);
	s_locks_lower_in(24,46) <= s_locks_lower_out(25,46);

		normal_cell_24_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,47),
			fetch              => s_fetch(24,47),
			data_in            => s_data_in(24,47),
			data_out           => s_data_out(24,47),
			out1               => s_out1(24,47),
			out2               => s_out2(24,47),
			lock_lower_row_out => s_locks_lower_out(24,47),
			lock_lower_row_in  => s_locks_lower_in(24,47),
			in1                => s_in1(24,47),
			in2                => s_in2(24,47),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(47)
		);
	s_in1(24,47)            <= s_out1(25,47);
	s_in2(24,47)            <= s_out2(25,48);
	s_locks_lower_in(24,47) <= s_locks_lower_out(25,47);

		normal_cell_24_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,48),
			fetch              => s_fetch(24,48),
			data_in            => s_data_in(24,48),
			data_out           => s_data_out(24,48),
			out1               => s_out1(24,48),
			out2               => s_out2(24,48),
			lock_lower_row_out => s_locks_lower_out(24,48),
			lock_lower_row_in  => s_locks_lower_in(24,48),
			in1                => s_in1(24,48),
			in2                => s_in2(24,48),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(48)
		);
	s_in1(24,48)            <= s_out1(25,48);
	s_in2(24,48)            <= s_out2(25,49);
	s_locks_lower_in(24,48) <= s_locks_lower_out(25,48);

		normal_cell_24_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,49),
			fetch              => s_fetch(24,49),
			data_in            => s_data_in(24,49),
			data_out           => s_data_out(24,49),
			out1               => s_out1(24,49),
			out2               => s_out2(24,49),
			lock_lower_row_out => s_locks_lower_out(24,49),
			lock_lower_row_in  => s_locks_lower_in(24,49),
			in1                => s_in1(24,49),
			in2                => s_in2(24,49),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(49)
		);
	s_in1(24,49)            <= s_out1(25,49);
	s_in2(24,49)            <= s_out2(25,50);
	s_locks_lower_in(24,49) <= s_locks_lower_out(25,49);

		normal_cell_24_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,50),
			fetch              => s_fetch(24,50),
			data_in            => s_data_in(24,50),
			data_out           => s_data_out(24,50),
			out1               => s_out1(24,50),
			out2               => s_out2(24,50),
			lock_lower_row_out => s_locks_lower_out(24,50),
			lock_lower_row_in  => s_locks_lower_in(24,50),
			in1                => s_in1(24,50),
			in2                => s_in2(24,50),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(50)
		);
	s_in1(24,50)            <= s_out1(25,50);
	s_in2(24,50)            <= s_out2(25,51);
	s_locks_lower_in(24,50) <= s_locks_lower_out(25,50);

		normal_cell_24_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,51),
			fetch              => s_fetch(24,51),
			data_in            => s_data_in(24,51),
			data_out           => s_data_out(24,51),
			out1               => s_out1(24,51),
			out2               => s_out2(24,51),
			lock_lower_row_out => s_locks_lower_out(24,51),
			lock_lower_row_in  => s_locks_lower_in(24,51),
			in1                => s_in1(24,51),
			in2                => s_in2(24,51),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(51)
		);
	s_in1(24,51)            <= s_out1(25,51);
	s_in2(24,51)            <= s_out2(25,52);
	s_locks_lower_in(24,51) <= s_locks_lower_out(25,51);

		normal_cell_24_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,52),
			fetch              => s_fetch(24,52),
			data_in            => s_data_in(24,52),
			data_out           => s_data_out(24,52),
			out1               => s_out1(24,52),
			out2               => s_out2(24,52),
			lock_lower_row_out => s_locks_lower_out(24,52),
			lock_lower_row_in  => s_locks_lower_in(24,52),
			in1                => s_in1(24,52),
			in2                => s_in2(24,52),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(52)
		);
	s_in1(24,52)            <= s_out1(25,52);
	s_in2(24,52)            <= s_out2(25,53);
	s_locks_lower_in(24,52) <= s_locks_lower_out(25,52);

		normal_cell_24_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,53),
			fetch              => s_fetch(24,53),
			data_in            => s_data_in(24,53),
			data_out           => s_data_out(24,53),
			out1               => s_out1(24,53),
			out2               => s_out2(24,53),
			lock_lower_row_out => s_locks_lower_out(24,53),
			lock_lower_row_in  => s_locks_lower_in(24,53),
			in1                => s_in1(24,53),
			in2                => s_in2(24,53),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(53)
		);
	s_in1(24,53)            <= s_out1(25,53);
	s_in2(24,53)            <= s_out2(25,54);
	s_locks_lower_in(24,53) <= s_locks_lower_out(25,53);

		normal_cell_24_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,54),
			fetch              => s_fetch(24,54),
			data_in            => s_data_in(24,54),
			data_out           => s_data_out(24,54),
			out1               => s_out1(24,54),
			out2               => s_out2(24,54),
			lock_lower_row_out => s_locks_lower_out(24,54),
			lock_lower_row_in  => s_locks_lower_in(24,54),
			in1                => s_in1(24,54),
			in2                => s_in2(24,54),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(54)
		);
	s_in1(24,54)            <= s_out1(25,54);
	s_in2(24,54)            <= s_out2(25,55);
	s_locks_lower_in(24,54) <= s_locks_lower_out(25,54);

		normal_cell_24_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,55),
			fetch              => s_fetch(24,55),
			data_in            => s_data_in(24,55),
			data_out           => s_data_out(24,55),
			out1               => s_out1(24,55),
			out2               => s_out2(24,55),
			lock_lower_row_out => s_locks_lower_out(24,55),
			lock_lower_row_in  => s_locks_lower_in(24,55),
			in1                => s_in1(24,55),
			in2                => s_in2(24,55),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(55)
		);
	s_in1(24,55)            <= s_out1(25,55);
	s_in2(24,55)            <= s_out2(25,56);
	s_locks_lower_in(24,55) <= s_locks_lower_out(25,55);

		normal_cell_24_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,56),
			fetch              => s_fetch(24,56),
			data_in            => s_data_in(24,56),
			data_out           => s_data_out(24,56),
			out1               => s_out1(24,56),
			out2               => s_out2(24,56),
			lock_lower_row_out => s_locks_lower_out(24,56),
			lock_lower_row_in  => s_locks_lower_in(24,56),
			in1                => s_in1(24,56),
			in2                => s_in2(24,56),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(56)
		);
	s_in1(24,56)            <= s_out1(25,56);
	s_in2(24,56)            <= s_out2(25,57);
	s_locks_lower_in(24,56) <= s_locks_lower_out(25,56);

		normal_cell_24_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,57),
			fetch              => s_fetch(24,57),
			data_in            => s_data_in(24,57),
			data_out           => s_data_out(24,57),
			out1               => s_out1(24,57),
			out2               => s_out2(24,57),
			lock_lower_row_out => s_locks_lower_out(24,57),
			lock_lower_row_in  => s_locks_lower_in(24,57),
			in1                => s_in1(24,57),
			in2                => s_in2(24,57),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(57)
		);
	s_in1(24,57)            <= s_out1(25,57);
	s_in2(24,57)            <= s_out2(25,58);
	s_locks_lower_in(24,57) <= s_locks_lower_out(25,57);

		normal_cell_24_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,58),
			fetch              => s_fetch(24,58),
			data_in            => s_data_in(24,58),
			data_out           => s_data_out(24,58),
			out1               => s_out1(24,58),
			out2               => s_out2(24,58),
			lock_lower_row_out => s_locks_lower_out(24,58),
			lock_lower_row_in  => s_locks_lower_in(24,58),
			in1                => s_in1(24,58),
			in2                => s_in2(24,58),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(58)
		);
	s_in1(24,58)            <= s_out1(25,58);
	s_in2(24,58)            <= s_out2(25,59);
	s_locks_lower_in(24,58) <= s_locks_lower_out(25,58);

		normal_cell_24_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,59),
			fetch              => s_fetch(24,59),
			data_in            => s_data_in(24,59),
			data_out           => s_data_out(24,59),
			out1               => s_out1(24,59),
			out2               => s_out2(24,59),
			lock_lower_row_out => s_locks_lower_out(24,59),
			lock_lower_row_in  => s_locks_lower_in(24,59),
			in1                => s_in1(24,59),
			in2                => s_in2(24,59),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(59)
		);
	s_in1(24,59)            <= s_out1(25,59);
	s_in2(24,59)            <= s_out2(25,60);
	s_locks_lower_in(24,59) <= s_locks_lower_out(25,59);

		last_col_cell_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(24,60),
			fetch              => s_fetch(24,60),
			data_in            => s_data_in(24,60),
			data_out           => s_data_out(24,60),
			out1               => s_out1(24,60),
			out2               => s_out2(24,60),
			lock_lower_row_out => s_locks_lower_out(24,60),
			lock_lower_row_in  => s_locks_lower_in(24,60),
			in1                => s_in1(24,60),
			in2                => (others => '0'),
			lock_row           => s_locks(24),
			piv_found          => s_piv_found,
			row_data           => s_row_data(24),
			col_data           => s_col_data(60)
		);
	s_in1(24,60)            <= s_out1(25,60);
	s_locks_lower_in(24,60) <= s_locks_lower_out(25,60);

		normal_cell_25_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,1),
			fetch              => s_fetch(25,1),
			data_in            => s_data_in(25,1),
			data_out           => s_data_out(25,1),
			out1               => s_out1(25,1),
			out2               => s_out2(25,1),
			lock_lower_row_out => s_locks_lower_out(25,1),
			lock_lower_row_in  => s_locks_lower_in(25,1),
			in1                => s_in1(25,1),
			in2                => s_in2(25,1),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(1)
		);
	s_in1(25,1)            <= s_out1(26,1);
	s_in2(25,1)            <= s_out2(26,2);
	s_locks_lower_in(25,1) <= s_locks_lower_out(26,1);

		normal_cell_25_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,2),
			fetch              => s_fetch(25,2),
			data_in            => s_data_in(25,2),
			data_out           => s_data_out(25,2),
			out1               => s_out1(25,2),
			out2               => s_out2(25,2),
			lock_lower_row_out => s_locks_lower_out(25,2),
			lock_lower_row_in  => s_locks_lower_in(25,2),
			in1                => s_in1(25,2),
			in2                => s_in2(25,2),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(2)
		);
	s_in1(25,2)            <= s_out1(26,2);
	s_in2(25,2)            <= s_out2(26,3);
	s_locks_lower_in(25,2) <= s_locks_lower_out(26,2);

		normal_cell_25_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,3),
			fetch              => s_fetch(25,3),
			data_in            => s_data_in(25,3),
			data_out           => s_data_out(25,3),
			out1               => s_out1(25,3),
			out2               => s_out2(25,3),
			lock_lower_row_out => s_locks_lower_out(25,3),
			lock_lower_row_in  => s_locks_lower_in(25,3),
			in1                => s_in1(25,3),
			in2                => s_in2(25,3),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(3)
		);
	s_in1(25,3)            <= s_out1(26,3);
	s_in2(25,3)            <= s_out2(26,4);
	s_locks_lower_in(25,3) <= s_locks_lower_out(26,3);

		normal_cell_25_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,4),
			fetch              => s_fetch(25,4),
			data_in            => s_data_in(25,4),
			data_out           => s_data_out(25,4),
			out1               => s_out1(25,4),
			out2               => s_out2(25,4),
			lock_lower_row_out => s_locks_lower_out(25,4),
			lock_lower_row_in  => s_locks_lower_in(25,4),
			in1                => s_in1(25,4),
			in2                => s_in2(25,4),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(4)
		);
	s_in1(25,4)            <= s_out1(26,4);
	s_in2(25,4)            <= s_out2(26,5);
	s_locks_lower_in(25,4) <= s_locks_lower_out(26,4);

		normal_cell_25_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,5),
			fetch              => s_fetch(25,5),
			data_in            => s_data_in(25,5),
			data_out           => s_data_out(25,5),
			out1               => s_out1(25,5),
			out2               => s_out2(25,5),
			lock_lower_row_out => s_locks_lower_out(25,5),
			lock_lower_row_in  => s_locks_lower_in(25,5),
			in1                => s_in1(25,5),
			in2                => s_in2(25,5),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(5)
		);
	s_in1(25,5)            <= s_out1(26,5);
	s_in2(25,5)            <= s_out2(26,6);
	s_locks_lower_in(25,5) <= s_locks_lower_out(26,5);

		normal_cell_25_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,6),
			fetch              => s_fetch(25,6),
			data_in            => s_data_in(25,6),
			data_out           => s_data_out(25,6),
			out1               => s_out1(25,6),
			out2               => s_out2(25,6),
			lock_lower_row_out => s_locks_lower_out(25,6),
			lock_lower_row_in  => s_locks_lower_in(25,6),
			in1                => s_in1(25,6),
			in2                => s_in2(25,6),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(6)
		);
	s_in1(25,6)            <= s_out1(26,6);
	s_in2(25,6)            <= s_out2(26,7);
	s_locks_lower_in(25,6) <= s_locks_lower_out(26,6);

		normal_cell_25_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,7),
			fetch              => s_fetch(25,7),
			data_in            => s_data_in(25,7),
			data_out           => s_data_out(25,7),
			out1               => s_out1(25,7),
			out2               => s_out2(25,7),
			lock_lower_row_out => s_locks_lower_out(25,7),
			lock_lower_row_in  => s_locks_lower_in(25,7),
			in1                => s_in1(25,7),
			in2                => s_in2(25,7),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(7)
		);
	s_in1(25,7)            <= s_out1(26,7);
	s_in2(25,7)            <= s_out2(26,8);
	s_locks_lower_in(25,7) <= s_locks_lower_out(26,7);

		normal_cell_25_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,8),
			fetch              => s_fetch(25,8),
			data_in            => s_data_in(25,8),
			data_out           => s_data_out(25,8),
			out1               => s_out1(25,8),
			out2               => s_out2(25,8),
			lock_lower_row_out => s_locks_lower_out(25,8),
			lock_lower_row_in  => s_locks_lower_in(25,8),
			in1                => s_in1(25,8),
			in2                => s_in2(25,8),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(8)
		);
	s_in1(25,8)            <= s_out1(26,8);
	s_in2(25,8)            <= s_out2(26,9);
	s_locks_lower_in(25,8) <= s_locks_lower_out(26,8);

		normal_cell_25_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,9),
			fetch              => s_fetch(25,9),
			data_in            => s_data_in(25,9),
			data_out           => s_data_out(25,9),
			out1               => s_out1(25,9),
			out2               => s_out2(25,9),
			lock_lower_row_out => s_locks_lower_out(25,9),
			lock_lower_row_in  => s_locks_lower_in(25,9),
			in1                => s_in1(25,9),
			in2                => s_in2(25,9),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(9)
		);
	s_in1(25,9)            <= s_out1(26,9);
	s_in2(25,9)            <= s_out2(26,10);
	s_locks_lower_in(25,9) <= s_locks_lower_out(26,9);

		normal_cell_25_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,10),
			fetch              => s_fetch(25,10),
			data_in            => s_data_in(25,10),
			data_out           => s_data_out(25,10),
			out1               => s_out1(25,10),
			out2               => s_out2(25,10),
			lock_lower_row_out => s_locks_lower_out(25,10),
			lock_lower_row_in  => s_locks_lower_in(25,10),
			in1                => s_in1(25,10),
			in2                => s_in2(25,10),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(10)
		);
	s_in1(25,10)            <= s_out1(26,10);
	s_in2(25,10)            <= s_out2(26,11);
	s_locks_lower_in(25,10) <= s_locks_lower_out(26,10);

		normal_cell_25_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,11),
			fetch              => s_fetch(25,11),
			data_in            => s_data_in(25,11),
			data_out           => s_data_out(25,11),
			out1               => s_out1(25,11),
			out2               => s_out2(25,11),
			lock_lower_row_out => s_locks_lower_out(25,11),
			lock_lower_row_in  => s_locks_lower_in(25,11),
			in1                => s_in1(25,11),
			in2                => s_in2(25,11),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(11)
		);
	s_in1(25,11)            <= s_out1(26,11);
	s_in2(25,11)            <= s_out2(26,12);
	s_locks_lower_in(25,11) <= s_locks_lower_out(26,11);

		normal_cell_25_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,12),
			fetch              => s_fetch(25,12),
			data_in            => s_data_in(25,12),
			data_out           => s_data_out(25,12),
			out1               => s_out1(25,12),
			out2               => s_out2(25,12),
			lock_lower_row_out => s_locks_lower_out(25,12),
			lock_lower_row_in  => s_locks_lower_in(25,12),
			in1                => s_in1(25,12),
			in2                => s_in2(25,12),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(12)
		);
	s_in1(25,12)            <= s_out1(26,12);
	s_in2(25,12)            <= s_out2(26,13);
	s_locks_lower_in(25,12) <= s_locks_lower_out(26,12);

		normal_cell_25_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,13),
			fetch              => s_fetch(25,13),
			data_in            => s_data_in(25,13),
			data_out           => s_data_out(25,13),
			out1               => s_out1(25,13),
			out2               => s_out2(25,13),
			lock_lower_row_out => s_locks_lower_out(25,13),
			lock_lower_row_in  => s_locks_lower_in(25,13),
			in1                => s_in1(25,13),
			in2                => s_in2(25,13),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(13)
		);
	s_in1(25,13)            <= s_out1(26,13);
	s_in2(25,13)            <= s_out2(26,14);
	s_locks_lower_in(25,13) <= s_locks_lower_out(26,13);

		normal_cell_25_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,14),
			fetch              => s_fetch(25,14),
			data_in            => s_data_in(25,14),
			data_out           => s_data_out(25,14),
			out1               => s_out1(25,14),
			out2               => s_out2(25,14),
			lock_lower_row_out => s_locks_lower_out(25,14),
			lock_lower_row_in  => s_locks_lower_in(25,14),
			in1                => s_in1(25,14),
			in2                => s_in2(25,14),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(14)
		);
	s_in1(25,14)            <= s_out1(26,14);
	s_in2(25,14)            <= s_out2(26,15);
	s_locks_lower_in(25,14) <= s_locks_lower_out(26,14);

		normal_cell_25_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,15),
			fetch              => s_fetch(25,15),
			data_in            => s_data_in(25,15),
			data_out           => s_data_out(25,15),
			out1               => s_out1(25,15),
			out2               => s_out2(25,15),
			lock_lower_row_out => s_locks_lower_out(25,15),
			lock_lower_row_in  => s_locks_lower_in(25,15),
			in1                => s_in1(25,15),
			in2                => s_in2(25,15),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(15)
		);
	s_in1(25,15)            <= s_out1(26,15);
	s_in2(25,15)            <= s_out2(26,16);
	s_locks_lower_in(25,15) <= s_locks_lower_out(26,15);

		normal_cell_25_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,16),
			fetch              => s_fetch(25,16),
			data_in            => s_data_in(25,16),
			data_out           => s_data_out(25,16),
			out1               => s_out1(25,16),
			out2               => s_out2(25,16),
			lock_lower_row_out => s_locks_lower_out(25,16),
			lock_lower_row_in  => s_locks_lower_in(25,16),
			in1                => s_in1(25,16),
			in2                => s_in2(25,16),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(16)
		);
	s_in1(25,16)            <= s_out1(26,16);
	s_in2(25,16)            <= s_out2(26,17);
	s_locks_lower_in(25,16) <= s_locks_lower_out(26,16);

		normal_cell_25_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,17),
			fetch              => s_fetch(25,17),
			data_in            => s_data_in(25,17),
			data_out           => s_data_out(25,17),
			out1               => s_out1(25,17),
			out2               => s_out2(25,17),
			lock_lower_row_out => s_locks_lower_out(25,17),
			lock_lower_row_in  => s_locks_lower_in(25,17),
			in1                => s_in1(25,17),
			in2                => s_in2(25,17),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(17)
		);
	s_in1(25,17)            <= s_out1(26,17);
	s_in2(25,17)            <= s_out2(26,18);
	s_locks_lower_in(25,17) <= s_locks_lower_out(26,17);

		normal_cell_25_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,18),
			fetch              => s_fetch(25,18),
			data_in            => s_data_in(25,18),
			data_out           => s_data_out(25,18),
			out1               => s_out1(25,18),
			out2               => s_out2(25,18),
			lock_lower_row_out => s_locks_lower_out(25,18),
			lock_lower_row_in  => s_locks_lower_in(25,18),
			in1                => s_in1(25,18),
			in2                => s_in2(25,18),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(18)
		);
	s_in1(25,18)            <= s_out1(26,18);
	s_in2(25,18)            <= s_out2(26,19);
	s_locks_lower_in(25,18) <= s_locks_lower_out(26,18);

		normal_cell_25_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,19),
			fetch              => s_fetch(25,19),
			data_in            => s_data_in(25,19),
			data_out           => s_data_out(25,19),
			out1               => s_out1(25,19),
			out2               => s_out2(25,19),
			lock_lower_row_out => s_locks_lower_out(25,19),
			lock_lower_row_in  => s_locks_lower_in(25,19),
			in1                => s_in1(25,19),
			in2                => s_in2(25,19),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(19)
		);
	s_in1(25,19)            <= s_out1(26,19);
	s_in2(25,19)            <= s_out2(26,20);
	s_locks_lower_in(25,19) <= s_locks_lower_out(26,19);

		normal_cell_25_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,20),
			fetch              => s_fetch(25,20),
			data_in            => s_data_in(25,20),
			data_out           => s_data_out(25,20),
			out1               => s_out1(25,20),
			out2               => s_out2(25,20),
			lock_lower_row_out => s_locks_lower_out(25,20),
			lock_lower_row_in  => s_locks_lower_in(25,20),
			in1                => s_in1(25,20),
			in2                => s_in2(25,20),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(20)
		);
	s_in1(25,20)            <= s_out1(26,20);
	s_in2(25,20)            <= s_out2(26,21);
	s_locks_lower_in(25,20) <= s_locks_lower_out(26,20);

		normal_cell_25_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,21),
			fetch              => s_fetch(25,21),
			data_in            => s_data_in(25,21),
			data_out           => s_data_out(25,21),
			out1               => s_out1(25,21),
			out2               => s_out2(25,21),
			lock_lower_row_out => s_locks_lower_out(25,21),
			lock_lower_row_in  => s_locks_lower_in(25,21),
			in1                => s_in1(25,21),
			in2                => s_in2(25,21),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(21)
		);
	s_in1(25,21)            <= s_out1(26,21);
	s_in2(25,21)            <= s_out2(26,22);
	s_locks_lower_in(25,21) <= s_locks_lower_out(26,21);

		normal_cell_25_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,22),
			fetch              => s_fetch(25,22),
			data_in            => s_data_in(25,22),
			data_out           => s_data_out(25,22),
			out1               => s_out1(25,22),
			out2               => s_out2(25,22),
			lock_lower_row_out => s_locks_lower_out(25,22),
			lock_lower_row_in  => s_locks_lower_in(25,22),
			in1                => s_in1(25,22),
			in2                => s_in2(25,22),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(22)
		);
	s_in1(25,22)            <= s_out1(26,22);
	s_in2(25,22)            <= s_out2(26,23);
	s_locks_lower_in(25,22) <= s_locks_lower_out(26,22);

		normal_cell_25_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,23),
			fetch              => s_fetch(25,23),
			data_in            => s_data_in(25,23),
			data_out           => s_data_out(25,23),
			out1               => s_out1(25,23),
			out2               => s_out2(25,23),
			lock_lower_row_out => s_locks_lower_out(25,23),
			lock_lower_row_in  => s_locks_lower_in(25,23),
			in1                => s_in1(25,23),
			in2                => s_in2(25,23),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(23)
		);
	s_in1(25,23)            <= s_out1(26,23);
	s_in2(25,23)            <= s_out2(26,24);
	s_locks_lower_in(25,23) <= s_locks_lower_out(26,23);

		normal_cell_25_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,24),
			fetch              => s_fetch(25,24),
			data_in            => s_data_in(25,24),
			data_out           => s_data_out(25,24),
			out1               => s_out1(25,24),
			out2               => s_out2(25,24),
			lock_lower_row_out => s_locks_lower_out(25,24),
			lock_lower_row_in  => s_locks_lower_in(25,24),
			in1                => s_in1(25,24),
			in2                => s_in2(25,24),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(24)
		);
	s_in1(25,24)            <= s_out1(26,24);
	s_in2(25,24)            <= s_out2(26,25);
	s_locks_lower_in(25,24) <= s_locks_lower_out(26,24);

		normal_cell_25_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,25),
			fetch              => s_fetch(25,25),
			data_in            => s_data_in(25,25),
			data_out           => s_data_out(25,25),
			out1               => s_out1(25,25),
			out2               => s_out2(25,25),
			lock_lower_row_out => s_locks_lower_out(25,25),
			lock_lower_row_in  => s_locks_lower_in(25,25),
			in1                => s_in1(25,25),
			in2                => s_in2(25,25),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(25)
		);
	s_in1(25,25)            <= s_out1(26,25);
	s_in2(25,25)            <= s_out2(26,26);
	s_locks_lower_in(25,25) <= s_locks_lower_out(26,25);

		normal_cell_25_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,26),
			fetch              => s_fetch(25,26),
			data_in            => s_data_in(25,26),
			data_out           => s_data_out(25,26),
			out1               => s_out1(25,26),
			out2               => s_out2(25,26),
			lock_lower_row_out => s_locks_lower_out(25,26),
			lock_lower_row_in  => s_locks_lower_in(25,26),
			in1                => s_in1(25,26),
			in2                => s_in2(25,26),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(26)
		);
	s_in1(25,26)            <= s_out1(26,26);
	s_in2(25,26)            <= s_out2(26,27);
	s_locks_lower_in(25,26) <= s_locks_lower_out(26,26);

		normal_cell_25_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,27),
			fetch              => s_fetch(25,27),
			data_in            => s_data_in(25,27),
			data_out           => s_data_out(25,27),
			out1               => s_out1(25,27),
			out2               => s_out2(25,27),
			lock_lower_row_out => s_locks_lower_out(25,27),
			lock_lower_row_in  => s_locks_lower_in(25,27),
			in1                => s_in1(25,27),
			in2                => s_in2(25,27),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(27)
		);
	s_in1(25,27)            <= s_out1(26,27);
	s_in2(25,27)            <= s_out2(26,28);
	s_locks_lower_in(25,27) <= s_locks_lower_out(26,27);

		normal_cell_25_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,28),
			fetch              => s_fetch(25,28),
			data_in            => s_data_in(25,28),
			data_out           => s_data_out(25,28),
			out1               => s_out1(25,28),
			out2               => s_out2(25,28),
			lock_lower_row_out => s_locks_lower_out(25,28),
			lock_lower_row_in  => s_locks_lower_in(25,28),
			in1                => s_in1(25,28),
			in2                => s_in2(25,28),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(28)
		);
	s_in1(25,28)            <= s_out1(26,28);
	s_in2(25,28)            <= s_out2(26,29);
	s_locks_lower_in(25,28) <= s_locks_lower_out(26,28);

		normal_cell_25_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,29),
			fetch              => s_fetch(25,29),
			data_in            => s_data_in(25,29),
			data_out           => s_data_out(25,29),
			out1               => s_out1(25,29),
			out2               => s_out2(25,29),
			lock_lower_row_out => s_locks_lower_out(25,29),
			lock_lower_row_in  => s_locks_lower_in(25,29),
			in1                => s_in1(25,29),
			in2                => s_in2(25,29),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(29)
		);
	s_in1(25,29)            <= s_out1(26,29);
	s_in2(25,29)            <= s_out2(26,30);
	s_locks_lower_in(25,29) <= s_locks_lower_out(26,29);

		normal_cell_25_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,30),
			fetch              => s_fetch(25,30),
			data_in            => s_data_in(25,30),
			data_out           => s_data_out(25,30),
			out1               => s_out1(25,30),
			out2               => s_out2(25,30),
			lock_lower_row_out => s_locks_lower_out(25,30),
			lock_lower_row_in  => s_locks_lower_in(25,30),
			in1                => s_in1(25,30),
			in2                => s_in2(25,30),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(30)
		);
	s_in1(25,30)            <= s_out1(26,30);
	s_in2(25,30)            <= s_out2(26,31);
	s_locks_lower_in(25,30) <= s_locks_lower_out(26,30);

		normal_cell_25_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,31),
			fetch              => s_fetch(25,31),
			data_in            => s_data_in(25,31),
			data_out           => s_data_out(25,31),
			out1               => s_out1(25,31),
			out2               => s_out2(25,31),
			lock_lower_row_out => s_locks_lower_out(25,31),
			lock_lower_row_in  => s_locks_lower_in(25,31),
			in1                => s_in1(25,31),
			in2                => s_in2(25,31),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(31)
		);
	s_in1(25,31)            <= s_out1(26,31);
	s_in2(25,31)            <= s_out2(26,32);
	s_locks_lower_in(25,31) <= s_locks_lower_out(26,31);

		normal_cell_25_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,32),
			fetch              => s_fetch(25,32),
			data_in            => s_data_in(25,32),
			data_out           => s_data_out(25,32),
			out1               => s_out1(25,32),
			out2               => s_out2(25,32),
			lock_lower_row_out => s_locks_lower_out(25,32),
			lock_lower_row_in  => s_locks_lower_in(25,32),
			in1                => s_in1(25,32),
			in2                => s_in2(25,32),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(32)
		);
	s_in1(25,32)            <= s_out1(26,32);
	s_in2(25,32)            <= s_out2(26,33);
	s_locks_lower_in(25,32) <= s_locks_lower_out(26,32);

		normal_cell_25_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,33),
			fetch              => s_fetch(25,33),
			data_in            => s_data_in(25,33),
			data_out           => s_data_out(25,33),
			out1               => s_out1(25,33),
			out2               => s_out2(25,33),
			lock_lower_row_out => s_locks_lower_out(25,33),
			lock_lower_row_in  => s_locks_lower_in(25,33),
			in1                => s_in1(25,33),
			in2                => s_in2(25,33),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(33)
		);
	s_in1(25,33)            <= s_out1(26,33);
	s_in2(25,33)            <= s_out2(26,34);
	s_locks_lower_in(25,33) <= s_locks_lower_out(26,33);

		normal_cell_25_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,34),
			fetch              => s_fetch(25,34),
			data_in            => s_data_in(25,34),
			data_out           => s_data_out(25,34),
			out1               => s_out1(25,34),
			out2               => s_out2(25,34),
			lock_lower_row_out => s_locks_lower_out(25,34),
			lock_lower_row_in  => s_locks_lower_in(25,34),
			in1                => s_in1(25,34),
			in2                => s_in2(25,34),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(34)
		);
	s_in1(25,34)            <= s_out1(26,34);
	s_in2(25,34)            <= s_out2(26,35);
	s_locks_lower_in(25,34) <= s_locks_lower_out(26,34);

		normal_cell_25_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,35),
			fetch              => s_fetch(25,35),
			data_in            => s_data_in(25,35),
			data_out           => s_data_out(25,35),
			out1               => s_out1(25,35),
			out2               => s_out2(25,35),
			lock_lower_row_out => s_locks_lower_out(25,35),
			lock_lower_row_in  => s_locks_lower_in(25,35),
			in1                => s_in1(25,35),
			in2                => s_in2(25,35),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(35)
		);
	s_in1(25,35)            <= s_out1(26,35);
	s_in2(25,35)            <= s_out2(26,36);
	s_locks_lower_in(25,35) <= s_locks_lower_out(26,35);

		normal_cell_25_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,36),
			fetch              => s_fetch(25,36),
			data_in            => s_data_in(25,36),
			data_out           => s_data_out(25,36),
			out1               => s_out1(25,36),
			out2               => s_out2(25,36),
			lock_lower_row_out => s_locks_lower_out(25,36),
			lock_lower_row_in  => s_locks_lower_in(25,36),
			in1                => s_in1(25,36),
			in2                => s_in2(25,36),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(36)
		);
	s_in1(25,36)            <= s_out1(26,36);
	s_in2(25,36)            <= s_out2(26,37);
	s_locks_lower_in(25,36) <= s_locks_lower_out(26,36);

		normal_cell_25_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,37),
			fetch              => s_fetch(25,37),
			data_in            => s_data_in(25,37),
			data_out           => s_data_out(25,37),
			out1               => s_out1(25,37),
			out2               => s_out2(25,37),
			lock_lower_row_out => s_locks_lower_out(25,37),
			lock_lower_row_in  => s_locks_lower_in(25,37),
			in1                => s_in1(25,37),
			in2                => s_in2(25,37),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(37)
		);
	s_in1(25,37)            <= s_out1(26,37);
	s_in2(25,37)            <= s_out2(26,38);
	s_locks_lower_in(25,37) <= s_locks_lower_out(26,37);

		normal_cell_25_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,38),
			fetch              => s_fetch(25,38),
			data_in            => s_data_in(25,38),
			data_out           => s_data_out(25,38),
			out1               => s_out1(25,38),
			out2               => s_out2(25,38),
			lock_lower_row_out => s_locks_lower_out(25,38),
			lock_lower_row_in  => s_locks_lower_in(25,38),
			in1                => s_in1(25,38),
			in2                => s_in2(25,38),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(38)
		);
	s_in1(25,38)            <= s_out1(26,38);
	s_in2(25,38)            <= s_out2(26,39);
	s_locks_lower_in(25,38) <= s_locks_lower_out(26,38);

		normal_cell_25_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,39),
			fetch              => s_fetch(25,39),
			data_in            => s_data_in(25,39),
			data_out           => s_data_out(25,39),
			out1               => s_out1(25,39),
			out2               => s_out2(25,39),
			lock_lower_row_out => s_locks_lower_out(25,39),
			lock_lower_row_in  => s_locks_lower_in(25,39),
			in1                => s_in1(25,39),
			in2                => s_in2(25,39),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(39)
		);
	s_in1(25,39)            <= s_out1(26,39);
	s_in2(25,39)            <= s_out2(26,40);
	s_locks_lower_in(25,39) <= s_locks_lower_out(26,39);

		normal_cell_25_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,40),
			fetch              => s_fetch(25,40),
			data_in            => s_data_in(25,40),
			data_out           => s_data_out(25,40),
			out1               => s_out1(25,40),
			out2               => s_out2(25,40),
			lock_lower_row_out => s_locks_lower_out(25,40),
			lock_lower_row_in  => s_locks_lower_in(25,40),
			in1                => s_in1(25,40),
			in2                => s_in2(25,40),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(40)
		);
	s_in1(25,40)            <= s_out1(26,40);
	s_in2(25,40)            <= s_out2(26,41);
	s_locks_lower_in(25,40) <= s_locks_lower_out(26,40);

		normal_cell_25_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,41),
			fetch              => s_fetch(25,41),
			data_in            => s_data_in(25,41),
			data_out           => s_data_out(25,41),
			out1               => s_out1(25,41),
			out2               => s_out2(25,41),
			lock_lower_row_out => s_locks_lower_out(25,41),
			lock_lower_row_in  => s_locks_lower_in(25,41),
			in1                => s_in1(25,41),
			in2                => s_in2(25,41),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(41)
		);
	s_in1(25,41)            <= s_out1(26,41);
	s_in2(25,41)            <= s_out2(26,42);
	s_locks_lower_in(25,41) <= s_locks_lower_out(26,41);

		normal_cell_25_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,42),
			fetch              => s_fetch(25,42),
			data_in            => s_data_in(25,42),
			data_out           => s_data_out(25,42),
			out1               => s_out1(25,42),
			out2               => s_out2(25,42),
			lock_lower_row_out => s_locks_lower_out(25,42),
			lock_lower_row_in  => s_locks_lower_in(25,42),
			in1                => s_in1(25,42),
			in2                => s_in2(25,42),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(42)
		);
	s_in1(25,42)            <= s_out1(26,42);
	s_in2(25,42)            <= s_out2(26,43);
	s_locks_lower_in(25,42) <= s_locks_lower_out(26,42);

		normal_cell_25_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,43),
			fetch              => s_fetch(25,43),
			data_in            => s_data_in(25,43),
			data_out           => s_data_out(25,43),
			out1               => s_out1(25,43),
			out2               => s_out2(25,43),
			lock_lower_row_out => s_locks_lower_out(25,43),
			lock_lower_row_in  => s_locks_lower_in(25,43),
			in1                => s_in1(25,43),
			in2                => s_in2(25,43),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(43)
		);
	s_in1(25,43)            <= s_out1(26,43);
	s_in2(25,43)            <= s_out2(26,44);
	s_locks_lower_in(25,43) <= s_locks_lower_out(26,43);

		normal_cell_25_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,44),
			fetch              => s_fetch(25,44),
			data_in            => s_data_in(25,44),
			data_out           => s_data_out(25,44),
			out1               => s_out1(25,44),
			out2               => s_out2(25,44),
			lock_lower_row_out => s_locks_lower_out(25,44),
			lock_lower_row_in  => s_locks_lower_in(25,44),
			in1                => s_in1(25,44),
			in2                => s_in2(25,44),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(44)
		);
	s_in1(25,44)            <= s_out1(26,44);
	s_in2(25,44)            <= s_out2(26,45);
	s_locks_lower_in(25,44) <= s_locks_lower_out(26,44);

		normal_cell_25_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,45),
			fetch              => s_fetch(25,45),
			data_in            => s_data_in(25,45),
			data_out           => s_data_out(25,45),
			out1               => s_out1(25,45),
			out2               => s_out2(25,45),
			lock_lower_row_out => s_locks_lower_out(25,45),
			lock_lower_row_in  => s_locks_lower_in(25,45),
			in1                => s_in1(25,45),
			in2                => s_in2(25,45),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(45)
		);
	s_in1(25,45)            <= s_out1(26,45);
	s_in2(25,45)            <= s_out2(26,46);
	s_locks_lower_in(25,45) <= s_locks_lower_out(26,45);

		normal_cell_25_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,46),
			fetch              => s_fetch(25,46),
			data_in            => s_data_in(25,46),
			data_out           => s_data_out(25,46),
			out1               => s_out1(25,46),
			out2               => s_out2(25,46),
			lock_lower_row_out => s_locks_lower_out(25,46),
			lock_lower_row_in  => s_locks_lower_in(25,46),
			in1                => s_in1(25,46),
			in2                => s_in2(25,46),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(46)
		);
	s_in1(25,46)            <= s_out1(26,46);
	s_in2(25,46)            <= s_out2(26,47);
	s_locks_lower_in(25,46) <= s_locks_lower_out(26,46);

		normal_cell_25_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,47),
			fetch              => s_fetch(25,47),
			data_in            => s_data_in(25,47),
			data_out           => s_data_out(25,47),
			out1               => s_out1(25,47),
			out2               => s_out2(25,47),
			lock_lower_row_out => s_locks_lower_out(25,47),
			lock_lower_row_in  => s_locks_lower_in(25,47),
			in1                => s_in1(25,47),
			in2                => s_in2(25,47),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(47)
		);
	s_in1(25,47)            <= s_out1(26,47);
	s_in2(25,47)            <= s_out2(26,48);
	s_locks_lower_in(25,47) <= s_locks_lower_out(26,47);

		normal_cell_25_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,48),
			fetch              => s_fetch(25,48),
			data_in            => s_data_in(25,48),
			data_out           => s_data_out(25,48),
			out1               => s_out1(25,48),
			out2               => s_out2(25,48),
			lock_lower_row_out => s_locks_lower_out(25,48),
			lock_lower_row_in  => s_locks_lower_in(25,48),
			in1                => s_in1(25,48),
			in2                => s_in2(25,48),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(48)
		);
	s_in1(25,48)            <= s_out1(26,48);
	s_in2(25,48)            <= s_out2(26,49);
	s_locks_lower_in(25,48) <= s_locks_lower_out(26,48);

		normal_cell_25_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,49),
			fetch              => s_fetch(25,49),
			data_in            => s_data_in(25,49),
			data_out           => s_data_out(25,49),
			out1               => s_out1(25,49),
			out2               => s_out2(25,49),
			lock_lower_row_out => s_locks_lower_out(25,49),
			lock_lower_row_in  => s_locks_lower_in(25,49),
			in1                => s_in1(25,49),
			in2                => s_in2(25,49),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(49)
		);
	s_in1(25,49)            <= s_out1(26,49);
	s_in2(25,49)            <= s_out2(26,50);
	s_locks_lower_in(25,49) <= s_locks_lower_out(26,49);

		normal_cell_25_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,50),
			fetch              => s_fetch(25,50),
			data_in            => s_data_in(25,50),
			data_out           => s_data_out(25,50),
			out1               => s_out1(25,50),
			out2               => s_out2(25,50),
			lock_lower_row_out => s_locks_lower_out(25,50),
			lock_lower_row_in  => s_locks_lower_in(25,50),
			in1                => s_in1(25,50),
			in2                => s_in2(25,50),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(50)
		);
	s_in1(25,50)            <= s_out1(26,50);
	s_in2(25,50)            <= s_out2(26,51);
	s_locks_lower_in(25,50) <= s_locks_lower_out(26,50);

		normal_cell_25_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,51),
			fetch              => s_fetch(25,51),
			data_in            => s_data_in(25,51),
			data_out           => s_data_out(25,51),
			out1               => s_out1(25,51),
			out2               => s_out2(25,51),
			lock_lower_row_out => s_locks_lower_out(25,51),
			lock_lower_row_in  => s_locks_lower_in(25,51),
			in1                => s_in1(25,51),
			in2                => s_in2(25,51),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(51)
		);
	s_in1(25,51)            <= s_out1(26,51);
	s_in2(25,51)            <= s_out2(26,52);
	s_locks_lower_in(25,51) <= s_locks_lower_out(26,51);

		normal_cell_25_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,52),
			fetch              => s_fetch(25,52),
			data_in            => s_data_in(25,52),
			data_out           => s_data_out(25,52),
			out1               => s_out1(25,52),
			out2               => s_out2(25,52),
			lock_lower_row_out => s_locks_lower_out(25,52),
			lock_lower_row_in  => s_locks_lower_in(25,52),
			in1                => s_in1(25,52),
			in2                => s_in2(25,52),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(52)
		);
	s_in1(25,52)            <= s_out1(26,52);
	s_in2(25,52)            <= s_out2(26,53);
	s_locks_lower_in(25,52) <= s_locks_lower_out(26,52);

		normal_cell_25_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,53),
			fetch              => s_fetch(25,53),
			data_in            => s_data_in(25,53),
			data_out           => s_data_out(25,53),
			out1               => s_out1(25,53),
			out2               => s_out2(25,53),
			lock_lower_row_out => s_locks_lower_out(25,53),
			lock_lower_row_in  => s_locks_lower_in(25,53),
			in1                => s_in1(25,53),
			in2                => s_in2(25,53),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(53)
		);
	s_in1(25,53)            <= s_out1(26,53);
	s_in2(25,53)            <= s_out2(26,54);
	s_locks_lower_in(25,53) <= s_locks_lower_out(26,53);

		normal_cell_25_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,54),
			fetch              => s_fetch(25,54),
			data_in            => s_data_in(25,54),
			data_out           => s_data_out(25,54),
			out1               => s_out1(25,54),
			out2               => s_out2(25,54),
			lock_lower_row_out => s_locks_lower_out(25,54),
			lock_lower_row_in  => s_locks_lower_in(25,54),
			in1                => s_in1(25,54),
			in2                => s_in2(25,54),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(54)
		);
	s_in1(25,54)            <= s_out1(26,54);
	s_in2(25,54)            <= s_out2(26,55);
	s_locks_lower_in(25,54) <= s_locks_lower_out(26,54);

		normal_cell_25_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,55),
			fetch              => s_fetch(25,55),
			data_in            => s_data_in(25,55),
			data_out           => s_data_out(25,55),
			out1               => s_out1(25,55),
			out2               => s_out2(25,55),
			lock_lower_row_out => s_locks_lower_out(25,55),
			lock_lower_row_in  => s_locks_lower_in(25,55),
			in1                => s_in1(25,55),
			in2                => s_in2(25,55),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(55)
		);
	s_in1(25,55)            <= s_out1(26,55);
	s_in2(25,55)            <= s_out2(26,56);
	s_locks_lower_in(25,55) <= s_locks_lower_out(26,55);

		normal_cell_25_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,56),
			fetch              => s_fetch(25,56),
			data_in            => s_data_in(25,56),
			data_out           => s_data_out(25,56),
			out1               => s_out1(25,56),
			out2               => s_out2(25,56),
			lock_lower_row_out => s_locks_lower_out(25,56),
			lock_lower_row_in  => s_locks_lower_in(25,56),
			in1                => s_in1(25,56),
			in2                => s_in2(25,56),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(56)
		);
	s_in1(25,56)            <= s_out1(26,56);
	s_in2(25,56)            <= s_out2(26,57);
	s_locks_lower_in(25,56) <= s_locks_lower_out(26,56);

		normal_cell_25_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,57),
			fetch              => s_fetch(25,57),
			data_in            => s_data_in(25,57),
			data_out           => s_data_out(25,57),
			out1               => s_out1(25,57),
			out2               => s_out2(25,57),
			lock_lower_row_out => s_locks_lower_out(25,57),
			lock_lower_row_in  => s_locks_lower_in(25,57),
			in1                => s_in1(25,57),
			in2                => s_in2(25,57),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(57)
		);
	s_in1(25,57)            <= s_out1(26,57);
	s_in2(25,57)            <= s_out2(26,58);
	s_locks_lower_in(25,57) <= s_locks_lower_out(26,57);

		normal_cell_25_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,58),
			fetch              => s_fetch(25,58),
			data_in            => s_data_in(25,58),
			data_out           => s_data_out(25,58),
			out1               => s_out1(25,58),
			out2               => s_out2(25,58),
			lock_lower_row_out => s_locks_lower_out(25,58),
			lock_lower_row_in  => s_locks_lower_in(25,58),
			in1                => s_in1(25,58),
			in2                => s_in2(25,58),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(58)
		);
	s_in1(25,58)            <= s_out1(26,58);
	s_in2(25,58)            <= s_out2(26,59);
	s_locks_lower_in(25,58) <= s_locks_lower_out(26,58);

		normal_cell_25_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,59),
			fetch              => s_fetch(25,59),
			data_in            => s_data_in(25,59),
			data_out           => s_data_out(25,59),
			out1               => s_out1(25,59),
			out2               => s_out2(25,59),
			lock_lower_row_out => s_locks_lower_out(25,59),
			lock_lower_row_in  => s_locks_lower_in(25,59),
			in1                => s_in1(25,59),
			in2                => s_in2(25,59),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(59)
		);
	s_in1(25,59)            <= s_out1(26,59);
	s_in2(25,59)            <= s_out2(26,60);
	s_locks_lower_in(25,59) <= s_locks_lower_out(26,59);

		last_col_cell_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(25,60),
			fetch              => s_fetch(25,60),
			data_in            => s_data_in(25,60),
			data_out           => s_data_out(25,60),
			out1               => s_out1(25,60),
			out2               => s_out2(25,60),
			lock_lower_row_out => s_locks_lower_out(25,60),
			lock_lower_row_in  => s_locks_lower_in(25,60),
			in1                => s_in1(25,60),
			in2                => (others => '0'),
			lock_row           => s_locks(25),
			piv_found          => s_piv_found,
			row_data           => s_row_data(25),
			col_data           => s_col_data(60)
		);
	s_in1(25,60)            <= s_out1(26,60);
	s_locks_lower_in(25,60) <= s_locks_lower_out(26,60);

		normal_cell_26_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,1),
			fetch              => s_fetch(26,1),
			data_in            => s_data_in(26,1),
			data_out           => s_data_out(26,1),
			out1               => s_out1(26,1),
			out2               => s_out2(26,1),
			lock_lower_row_out => s_locks_lower_out(26,1),
			lock_lower_row_in  => s_locks_lower_in(26,1),
			in1                => s_in1(26,1),
			in2                => s_in2(26,1),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(1)
		);
	s_in1(26,1)            <= s_out1(27,1);
	s_in2(26,1)            <= s_out2(27,2);
	s_locks_lower_in(26,1) <= s_locks_lower_out(27,1);

		normal_cell_26_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,2),
			fetch              => s_fetch(26,2),
			data_in            => s_data_in(26,2),
			data_out           => s_data_out(26,2),
			out1               => s_out1(26,2),
			out2               => s_out2(26,2),
			lock_lower_row_out => s_locks_lower_out(26,2),
			lock_lower_row_in  => s_locks_lower_in(26,2),
			in1                => s_in1(26,2),
			in2                => s_in2(26,2),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(2)
		);
	s_in1(26,2)            <= s_out1(27,2);
	s_in2(26,2)            <= s_out2(27,3);
	s_locks_lower_in(26,2) <= s_locks_lower_out(27,2);

		normal_cell_26_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,3),
			fetch              => s_fetch(26,3),
			data_in            => s_data_in(26,3),
			data_out           => s_data_out(26,3),
			out1               => s_out1(26,3),
			out2               => s_out2(26,3),
			lock_lower_row_out => s_locks_lower_out(26,3),
			lock_lower_row_in  => s_locks_lower_in(26,3),
			in1                => s_in1(26,3),
			in2                => s_in2(26,3),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(3)
		);
	s_in1(26,3)            <= s_out1(27,3);
	s_in2(26,3)            <= s_out2(27,4);
	s_locks_lower_in(26,3) <= s_locks_lower_out(27,3);

		normal_cell_26_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,4),
			fetch              => s_fetch(26,4),
			data_in            => s_data_in(26,4),
			data_out           => s_data_out(26,4),
			out1               => s_out1(26,4),
			out2               => s_out2(26,4),
			lock_lower_row_out => s_locks_lower_out(26,4),
			lock_lower_row_in  => s_locks_lower_in(26,4),
			in1                => s_in1(26,4),
			in2                => s_in2(26,4),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(4)
		);
	s_in1(26,4)            <= s_out1(27,4);
	s_in2(26,4)            <= s_out2(27,5);
	s_locks_lower_in(26,4) <= s_locks_lower_out(27,4);

		normal_cell_26_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,5),
			fetch              => s_fetch(26,5),
			data_in            => s_data_in(26,5),
			data_out           => s_data_out(26,5),
			out1               => s_out1(26,5),
			out2               => s_out2(26,5),
			lock_lower_row_out => s_locks_lower_out(26,5),
			lock_lower_row_in  => s_locks_lower_in(26,5),
			in1                => s_in1(26,5),
			in2                => s_in2(26,5),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(5)
		);
	s_in1(26,5)            <= s_out1(27,5);
	s_in2(26,5)            <= s_out2(27,6);
	s_locks_lower_in(26,5) <= s_locks_lower_out(27,5);

		normal_cell_26_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,6),
			fetch              => s_fetch(26,6),
			data_in            => s_data_in(26,6),
			data_out           => s_data_out(26,6),
			out1               => s_out1(26,6),
			out2               => s_out2(26,6),
			lock_lower_row_out => s_locks_lower_out(26,6),
			lock_lower_row_in  => s_locks_lower_in(26,6),
			in1                => s_in1(26,6),
			in2                => s_in2(26,6),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(6)
		);
	s_in1(26,6)            <= s_out1(27,6);
	s_in2(26,6)            <= s_out2(27,7);
	s_locks_lower_in(26,6) <= s_locks_lower_out(27,6);

		normal_cell_26_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,7),
			fetch              => s_fetch(26,7),
			data_in            => s_data_in(26,7),
			data_out           => s_data_out(26,7),
			out1               => s_out1(26,7),
			out2               => s_out2(26,7),
			lock_lower_row_out => s_locks_lower_out(26,7),
			lock_lower_row_in  => s_locks_lower_in(26,7),
			in1                => s_in1(26,7),
			in2                => s_in2(26,7),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(7)
		);
	s_in1(26,7)            <= s_out1(27,7);
	s_in2(26,7)            <= s_out2(27,8);
	s_locks_lower_in(26,7) <= s_locks_lower_out(27,7);

		normal_cell_26_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,8),
			fetch              => s_fetch(26,8),
			data_in            => s_data_in(26,8),
			data_out           => s_data_out(26,8),
			out1               => s_out1(26,8),
			out2               => s_out2(26,8),
			lock_lower_row_out => s_locks_lower_out(26,8),
			lock_lower_row_in  => s_locks_lower_in(26,8),
			in1                => s_in1(26,8),
			in2                => s_in2(26,8),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(8)
		);
	s_in1(26,8)            <= s_out1(27,8);
	s_in2(26,8)            <= s_out2(27,9);
	s_locks_lower_in(26,8) <= s_locks_lower_out(27,8);

		normal_cell_26_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,9),
			fetch              => s_fetch(26,9),
			data_in            => s_data_in(26,9),
			data_out           => s_data_out(26,9),
			out1               => s_out1(26,9),
			out2               => s_out2(26,9),
			lock_lower_row_out => s_locks_lower_out(26,9),
			lock_lower_row_in  => s_locks_lower_in(26,9),
			in1                => s_in1(26,9),
			in2                => s_in2(26,9),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(9)
		);
	s_in1(26,9)            <= s_out1(27,9);
	s_in2(26,9)            <= s_out2(27,10);
	s_locks_lower_in(26,9) <= s_locks_lower_out(27,9);

		normal_cell_26_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,10),
			fetch              => s_fetch(26,10),
			data_in            => s_data_in(26,10),
			data_out           => s_data_out(26,10),
			out1               => s_out1(26,10),
			out2               => s_out2(26,10),
			lock_lower_row_out => s_locks_lower_out(26,10),
			lock_lower_row_in  => s_locks_lower_in(26,10),
			in1                => s_in1(26,10),
			in2                => s_in2(26,10),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(10)
		);
	s_in1(26,10)            <= s_out1(27,10);
	s_in2(26,10)            <= s_out2(27,11);
	s_locks_lower_in(26,10) <= s_locks_lower_out(27,10);

		normal_cell_26_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,11),
			fetch              => s_fetch(26,11),
			data_in            => s_data_in(26,11),
			data_out           => s_data_out(26,11),
			out1               => s_out1(26,11),
			out2               => s_out2(26,11),
			lock_lower_row_out => s_locks_lower_out(26,11),
			lock_lower_row_in  => s_locks_lower_in(26,11),
			in1                => s_in1(26,11),
			in2                => s_in2(26,11),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(11)
		);
	s_in1(26,11)            <= s_out1(27,11);
	s_in2(26,11)            <= s_out2(27,12);
	s_locks_lower_in(26,11) <= s_locks_lower_out(27,11);

		normal_cell_26_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,12),
			fetch              => s_fetch(26,12),
			data_in            => s_data_in(26,12),
			data_out           => s_data_out(26,12),
			out1               => s_out1(26,12),
			out2               => s_out2(26,12),
			lock_lower_row_out => s_locks_lower_out(26,12),
			lock_lower_row_in  => s_locks_lower_in(26,12),
			in1                => s_in1(26,12),
			in2                => s_in2(26,12),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(12)
		);
	s_in1(26,12)            <= s_out1(27,12);
	s_in2(26,12)            <= s_out2(27,13);
	s_locks_lower_in(26,12) <= s_locks_lower_out(27,12);

		normal_cell_26_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,13),
			fetch              => s_fetch(26,13),
			data_in            => s_data_in(26,13),
			data_out           => s_data_out(26,13),
			out1               => s_out1(26,13),
			out2               => s_out2(26,13),
			lock_lower_row_out => s_locks_lower_out(26,13),
			lock_lower_row_in  => s_locks_lower_in(26,13),
			in1                => s_in1(26,13),
			in2                => s_in2(26,13),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(13)
		);
	s_in1(26,13)            <= s_out1(27,13);
	s_in2(26,13)            <= s_out2(27,14);
	s_locks_lower_in(26,13) <= s_locks_lower_out(27,13);

		normal_cell_26_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,14),
			fetch              => s_fetch(26,14),
			data_in            => s_data_in(26,14),
			data_out           => s_data_out(26,14),
			out1               => s_out1(26,14),
			out2               => s_out2(26,14),
			lock_lower_row_out => s_locks_lower_out(26,14),
			lock_lower_row_in  => s_locks_lower_in(26,14),
			in1                => s_in1(26,14),
			in2                => s_in2(26,14),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(14)
		);
	s_in1(26,14)            <= s_out1(27,14);
	s_in2(26,14)            <= s_out2(27,15);
	s_locks_lower_in(26,14) <= s_locks_lower_out(27,14);

		normal_cell_26_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,15),
			fetch              => s_fetch(26,15),
			data_in            => s_data_in(26,15),
			data_out           => s_data_out(26,15),
			out1               => s_out1(26,15),
			out2               => s_out2(26,15),
			lock_lower_row_out => s_locks_lower_out(26,15),
			lock_lower_row_in  => s_locks_lower_in(26,15),
			in1                => s_in1(26,15),
			in2                => s_in2(26,15),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(15)
		);
	s_in1(26,15)            <= s_out1(27,15);
	s_in2(26,15)            <= s_out2(27,16);
	s_locks_lower_in(26,15) <= s_locks_lower_out(27,15);

		normal_cell_26_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,16),
			fetch              => s_fetch(26,16),
			data_in            => s_data_in(26,16),
			data_out           => s_data_out(26,16),
			out1               => s_out1(26,16),
			out2               => s_out2(26,16),
			lock_lower_row_out => s_locks_lower_out(26,16),
			lock_lower_row_in  => s_locks_lower_in(26,16),
			in1                => s_in1(26,16),
			in2                => s_in2(26,16),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(16)
		);
	s_in1(26,16)            <= s_out1(27,16);
	s_in2(26,16)            <= s_out2(27,17);
	s_locks_lower_in(26,16) <= s_locks_lower_out(27,16);

		normal_cell_26_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,17),
			fetch              => s_fetch(26,17),
			data_in            => s_data_in(26,17),
			data_out           => s_data_out(26,17),
			out1               => s_out1(26,17),
			out2               => s_out2(26,17),
			lock_lower_row_out => s_locks_lower_out(26,17),
			lock_lower_row_in  => s_locks_lower_in(26,17),
			in1                => s_in1(26,17),
			in2                => s_in2(26,17),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(17)
		);
	s_in1(26,17)            <= s_out1(27,17);
	s_in2(26,17)            <= s_out2(27,18);
	s_locks_lower_in(26,17) <= s_locks_lower_out(27,17);

		normal_cell_26_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,18),
			fetch              => s_fetch(26,18),
			data_in            => s_data_in(26,18),
			data_out           => s_data_out(26,18),
			out1               => s_out1(26,18),
			out2               => s_out2(26,18),
			lock_lower_row_out => s_locks_lower_out(26,18),
			lock_lower_row_in  => s_locks_lower_in(26,18),
			in1                => s_in1(26,18),
			in2                => s_in2(26,18),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(18)
		);
	s_in1(26,18)            <= s_out1(27,18);
	s_in2(26,18)            <= s_out2(27,19);
	s_locks_lower_in(26,18) <= s_locks_lower_out(27,18);

		normal_cell_26_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,19),
			fetch              => s_fetch(26,19),
			data_in            => s_data_in(26,19),
			data_out           => s_data_out(26,19),
			out1               => s_out1(26,19),
			out2               => s_out2(26,19),
			lock_lower_row_out => s_locks_lower_out(26,19),
			lock_lower_row_in  => s_locks_lower_in(26,19),
			in1                => s_in1(26,19),
			in2                => s_in2(26,19),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(19)
		);
	s_in1(26,19)            <= s_out1(27,19);
	s_in2(26,19)            <= s_out2(27,20);
	s_locks_lower_in(26,19) <= s_locks_lower_out(27,19);

		normal_cell_26_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,20),
			fetch              => s_fetch(26,20),
			data_in            => s_data_in(26,20),
			data_out           => s_data_out(26,20),
			out1               => s_out1(26,20),
			out2               => s_out2(26,20),
			lock_lower_row_out => s_locks_lower_out(26,20),
			lock_lower_row_in  => s_locks_lower_in(26,20),
			in1                => s_in1(26,20),
			in2                => s_in2(26,20),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(20)
		);
	s_in1(26,20)            <= s_out1(27,20);
	s_in2(26,20)            <= s_out2(27,21);
	s_locks_lower_in(26,20) <= s_locks_lower_out(27,20);

		normal_cell_26_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,21),
			fetch              => s_fetch(26,21),
			data_in            => s_data_in(26,21),
			data_out           => s_data_out(26,21),
			out1               => s_out1(26,21),
			out2               => s_out2(26,21),
			lock_lower_row_out => s_locks_lower_out(26,21),
			lock_lower_row_in  => s_locks_lower_in(26,21),
			in1                => s_in1(26,21),
			in2                => s_in2(26,21),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(21)
		);
	s_in1(26,21)            <= s_out1(27,21);
	s_in2(26,21)            <= s_out2(27,22);
	s_locks_lower_in(26,21) <= s_locks_lower_out(27,21);

		normal_cell_26_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,22),
			fetch              => s_fetch(26,22),
			data_in            => s_data_in(26,22),
			data_out           => s_data_out(26,22),
			out1               => s_out1(26,22),
			out2               => s_out2(26,22),
			lock_lower_row_out => s_locks_lower_out(26,22),
			lock_lower_row_in  => s_locks_lower_in(26,22),
			in1                => s_in1(26,22),
			in2                => s_in2(26,22),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(22)
		);
	s_in1(26,22)            <= s_out1(27,22);
	s_in2(26,22)            <= s_out2(27,23);
	s_locks_lower_in(26,22) <= s_locks_lower_out(27,22);

		normal_cell_26_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,23),
			fetch              => s_fetch(26,23),
			data_in            => s_data_in(26,23),
			data_out           => s_data_out(26,23),
			out1               => s_out1(26,23),
			out2               => s_out2(26,23),
			lock_lower_row_out => s_locks_lower_out(26,23),
			lock_lower_row_in  => s_locks_lower_in(26,23),
			in1                => s_in1(26,23),
			in2                => s_in2(26,23),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(23)
		);
	s_in1(26,23)            <= s_out1(27,23);
	s_in2(26,23)            <= s_out2(27,24);
	s_locks_lower_in(26,23) <= s_locks_lower_out(27,23);

		normal_cell_26_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,24),
			fetch              => s_fetch(26,24),
			data_in            => s_data_in(26,24),
			data_out           => s_data_out(26,24),
			out1               => s_out1(26,24),
			out2               => s_out2(26,24),
			lock_lower_row_out => s_locks_lower_out(26,24),
			lock_lower_row_in  => s_locks_lower_in(26,24),
			in1                => s_in1(26,24),
			in2                => s_in2(26,24),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(24)
		);
	s_in1(26,24)            <= s_out1(27,24);
	s_in2(26,24)            <= s_out2(27,25);
	s_locks_lower_in(26,24) <= s_locks_lower_out(27,24);

		normal_cell_26_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,25),
			fetch              => s_fetch(26,25),
			data_in            => s_data_in(26,25),
			data_out           => s_data_out(26,25),
			out1               => s_out1(26,25),
			out2               => s_out2(26,25),
			lock_lower_row_out => s_locks_lower_out(26,25),
			lock_lower_row_in  => s_locks_lower_in(26,25),
			in1                => s_in1(26,25),
			in2                => s_in2(26,25),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(25)
		);
	s_in1(26,25)            <= s_out1(27,25);
	s_in2(26,25)            <= s_out2(27,26);
	s_locks_lower_in(26,25) <= s_locks_lower_out(27,25);

		normal_cell_26_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,26),
			fetch              => s_fetch(26,26),
			data_in            => s_data_in(26,26),
			data_out           => s_data_out(26,26),
			out1               => s_out1(26,26),
			out2               => s_out2(26,26),
			lock_lower_row_out => s_locks_lower_out(26,26),
			lock_lower_row_in  => s_locks_lower_in(26,26),
			in1                => s_in1(26,26),
			in2                => s_in2(26,26),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(26)
		);
	s_in1(26,26)            <= s_out1(27,26);
	s_in2(26,26)            <= s_out2(27,27);
	s_locks_lower_in(26,26) <= s_locks_lower_out(27,26);

		normal_cell_26_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,27),
			fetch              => s_fetch(26,27),
			data_in            => s_data_in(26,27),
			data_out           => s_data_out(26,27),
			out1               => s_out1(26,27),
			out2               => s_out2(26,27),
			lock_lower_row_out => s_locks_lower_out(26,27),
			lock_lower_row_in  => s_locks_lower_in(26,27),
			in1                => s_in1(26,27),
			in2                => s_in2(26,27),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(27)
		);
	s_in1(26,27)            <= s_out1(27,27);
	s_in2(26,27)            <= s_out2(27,28);
	s_locks_lower_in(26,27) <= s_locks_lower_out(27,27);

		normal_cell_26_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,28),
			fetch              => s_fetch(26,28),
			data_in            => s_data_in(26,28),
			data_out           => s_data_out(26,28),
			out1               => s_out1(26,28),
			out2               => s_out2(26,28),
			lock_lower_row_out => s_locks_lower_out(26,28),
			lock_lower_row_in  => s_locks_lower_in(26,28),
			in1                => s_in1(26,28),
			in2                => s_in2(26,28),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(28)
		);
	s_in1(26,28)            <= s_out1(27,28);
	s_in2(26,28)            <= s_out2(27,29);
	s_locks_lower_in(26,28) <= s_locks_lower_out(27,28);

		normal_cell_26_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,29),
			fetch              => s_fetch(26,29),
			data_in            => s_data_in(26,29),
			data_out           => s_data_out(26,29),
			out1               => s_out1(26,29),
			out2               => s_out2(26,29),
			lock_lower_row_out => s_locks_lower_out(26,29),
			lock_lower_row_in  => s_locks_lower_in(26,29),
			in1                => s_in1(26,29),
			in2                => s_in2(26,29),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(29)
		);
	s_in1(26,29)            <= s_out1(27,29);
	s_in2(26,29)            <= s_out2(27,30);
	s_locks_lower_in(26,29) <= s_locks_lower_out(27,29);

		normal_cell_26_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,30),
			fetch              => s_fetch(26,30),
			data_in            => s_data_in(26,30),
			data_out           => s_data_out(26,30),
			out1               => s_out1(26,30),
			out2               => s_out2(26,30),
			lock_lower_row_out => s_locks_lower_out(26,30),
			lock_lower_row_in  => s_locks_lower_in(26,30),
			in1                => s_in1(26,30),
			in2                => s_in2(26,30),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(30)
		);
	s_in1(26,30)            <= s_out1(27,30);
	s_in2(26,30)            <= s_out2(27,31);
	s_locks_lower_in(26,30) <= s_locks_lower_out(27,30);

		normal_cell_26_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,31),
			fetch              => s_fetch(26,31),
			data_in            => s_data_in(26,31),
			data_out           => s_data_out(26,31),
			out1               => s_out1(26,31),
			out2               => s_out2(26,31),
			lock_lower_row_out => s_locks_lower_out(26,31),
			lock_lower_row_in  => s_locks_lower_in(26,31),
			in1                => s_in1(26,31),
			in2                => s_in2(26,31),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(31)
		);
	s_in1(26,31)            <= s_out1(27,31);
	s_in2(26,31)            <= s_out2(27,32);
	s_locks_lower_in(26,31) <= s_locks_lower_out(27,31);

		normal_cell_26_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,32),
			fetch              => s_fetch(26,32),
			data_in            => s_data_in(26,32),
			data_out           => s_data_out(26,32),
			out1               => s_out1(26,32),
			out2               => s_out2(26,32),
			lock_lower_row_out => s_locks_lower_out(26,32),
			lock_lower_row_in  => s_locks_lower_in(26,32),
			in1                => s_in1(26,32),
			in2                => s_in2(26,32),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(32)
		);
	s_in1(26,32)            <= s_out1(27,32);
	s_in2(26,32)            <= s_out2(27,33);
	s_locks_lower_in(26,32) <= s_locks_lower_out(27,32);

		normal_cell_26_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,33),
			fetch              => s_fetch(26,33),
			data_in            => s_data_in(26,33),
			data_out           => s_data_out(26,33),
			out1               => s_out1(26,33),
			out2               => s_out2(26,33),
			lock_lower_row_out => s_locks_lower_out(26,33),
			lock_lower_row_in  => s_locks_lower_in(26,33),
			in1                => s_in1(26,33),
			in2                => s_in2(26,33),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(33)
		);
	s_in1(26,33)            <= s_out1(27,33);
	s_in2(26,33)            <= s_out2(27,34);
	s_locks_lower_in(26,33) <= s_locks_lower_out(27,33);

		normal_cell_26_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,34),
			fetch              => s_fetch(26,34),
			data_in            => s_data_in(26,34),
			data_out           => s_data_out(26,34),
			out1               => s_out1(26,34),
			out2               => s_out2(26,34),
			lock_lower_row_out => s_locks_lower_out(26,34),
			lock_lower_row_in  => s_locks_lower_in(26,34),
			in1                => s_in1(26,34),
			in2                => s_in2(26,34),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(34)
		);
	s_in1(26,34)            <= s_out1(27,34);
	s_in2(26,34)            <= s_out2(27,35);
	s_locks_lower_in(26,34) <= s_locks_lower_out(27,34);

		normal_cell_26_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,35),
			fetch              => s_fetch(26,35),
			data_in            => s_data_in(26,35),
			data_out           => s_data_out(26,35),
			out1               => s_out1(26,35),
			out2               => s_out2(26,35),
			lock_lower_row_out => s_locks_lower_out(26,35),
			lock_lower_row_in  => s_locks_lower_in(26,35),
			in1                => s_in1(26,35),
			in2                => s_in2(26,35),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(35)
		);
	s_in1(26,35)            <= s_out1(27,35);
	s_in2(26,35)            <= s_out2(27,36);
	s_locks_lower_in(26,35) <= s_locks_lower_out(27,35);

		normal_cell_26_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,36),
			fetch              => s_fetch(26,36),
			data_in            => s_data_in(26,36),
			data_out           => s_data_out(26,36),
			out1               => s_out1(26,36),
			out2               => s_out2(26,36),
			lock_lower_row_out => s_locks_lower_out(26,36),
			lock_lower_row_in  => s_locks_lower_in(26,36),
			in1                => s_in1(26,36),
			in2                => s_in2(26,36),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(36)
		);
	s_in1(26,36)            <= s_out1(27,36);
	s_in2(26,36)            <= s_out2(27,37);
	s_locks_lower_in(26,36) <= s_locks_lower_out(27,36);

		normal_cell_26_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,37),
			fetch              => s_fetch(26,37),
			data_in            => s_data_in(26,37),
			data_out           => s_data_out(26,37),
			out1               => s_out1(26,37),
			out2               => s_out2(26,37),
			lock_lower_row_out => s_locks_lower_out(26,37),
			lock_lower_row_in  => s_locks_lower_in(26,37),
			in1                => s_in1(26,37),
			in2                => s_in2(26,37),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(37)
		);
	s_in1(26,37)            <= s_out1(27,37);
	s_in2(26,37)            <= s_out2(27,38);
	s_locks_lower_in(26,37) <= s_locks_lower_out(27,37);

		normal_cell_26_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,38),
			fetch              => s_fetch(26,38),
			data_in            => s_data_in(26,38),
			data_out           => s_data_out(26,38),
			out1               => s_out1(26,38),
			out2               => s_out2(26,38),
			lock_lower_row_out => s_locks_lower_out(26,38),
			lock_lower_row_in  => s_locks_lower_in(26,38),
			in1                => s_in1(26,38),
			in2                => s_in2(26,38),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(38)
		);
	s_in1(26,38)            <= s_out1(27,38);
	s_in2(26,38)            <= s_out2(27,39);
	s_locks_lower_in(26,38) <= s_locks_lower_out(27,38);

		normal_cell_26_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,39),
			fetch              => s_fetch(26,39),
			data_in            => s_data_in(26,39),
			data_out           => s_data_out(26,39),
			out1               => s_out1(26,39),
			out2               => s_out2(26,39),
			lock_lower_row_out => s_locks_lower_out(26,39),
			lock_lower_row_in  => s_locks_lower_in(26,39),
			in1                => s_in1(26,39),
			in2                => s_in2(26,39),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(39)
		);
	s_in1(26,39)            <= s_out1(27,39);
	s_in2(26,39)            <= s_out2(27,40);
	s_locks_lower_in(26,39) <= s_locks_lower_out(27,39);

		normal_cell_26_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,40),
			fetch              => s_fetch(26,40),
			data_in            => s_data_in(26,40),
			data_out           => s_data_out(26,40),
			out1               => s_out1(26,40),
			out2               => s_out2(26,40),
			lock_lower_row_out => s_locks_lower_out(26,40),
			lock_lower_row_in  => s_locks_lower_in(26,40),
			in1                => s_in1(26,40),
			in2                => s_in2(26,40),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(40)
		);
	s_in1(26,40)            <= s_out1(27,40);
	s_in2(26,40)            <= s_out2(27,41);
	s_locks_lower_in(26,40) <= s_locks_lower_out(27,40);

		normal_cell_26_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,41),
			fetch              => s_fetch(26,41),
			data_in            => s_data_in(26,41),
			data_out           => s_data_out(26,41),
			out1               => s_out1(26,41),
			out2               => s_out2(26,41),
			lock_lower_row_out => s_locks_lower_out(26,41),
			lock_lower_row_in  => s_locks_lower_in(26,41),
			in1                => s_in1(26,41),
			in2                => s_in2(26,41),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(41)
		);
	s_in1(26,41)            <= s_out1(27,41);
	s_in2(26,41)            <= s_out2(27,42);
	s_locks_lower_in(26,41) <= s_locks_lower_out(27,41);

		normal_cell_26_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,42),
			fetch              => s_fetch(26,42),
			data_in            => s_data_in(26,42),
			data_out           => s_data_out(26,42),
			out1               => s_out1(26,42),
			out2               => s_out2(26,42),
			lock_lower_row_out => s_locks_lower_out(26,42),
			lock_lower_row_in  => s_locks_lower_in(26,42),
			in1                => s_in1(26,42),
			in2                => s_in2(26,42),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(42)
		);
	s_in1(26,42)            <= s_out1(27,42);
	s_in2(26,42)            <= s_out2(27,43);
	s_locks_lower_in(26,42) <= s_locks_lower_out(27,42);

		normal_cell_26_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,43),
			fetch              => s_fetch(26,43),
			data_in            => s_data_in(26,43),
			data_out           => s_data_out(26,43),
			out1               => s_out1(26,43),
			out2               => s_out2(26,43),
			lock_lower_row_out => s_locks_lower_out(26,43),
			lock_lower_row_in  => s_locks_lower_in(26,43),
			in1                => s_in1(26,43),
			in2                => s_in2(26,43),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(43)
		);
	s_in1(26,43)            <= s_out1(27,43);
	s_in2(26,43)            <= s_out2(27,44);
	s_locks_lower_in(26,43) <= s_locks_lower_out(27,43);

		normal_cell_26_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,44),
			fetch              => s_fetch(26,44),
			data_in            => s_data_in(26,44),
			data_out           => s_data_out(26,44),
			out1               => s_out1(26,44),
			out2               => s_out2(26,44),
			lock_lower_row_out => s_locks_lower_out(26,44),
			lock_lower_row_in  => s_locks_lower_in(26,44),
			in1                => s_in1(26,44),
			in2                => s_in2(26,44),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(44)
		);
	s_in1(26,44)            <= s_out1(27,44);
	s_in2(26,44)            <= s_out2(27,45);
	s_locks_lower_in(26,44) <= s_locks_lower_out(27,44);

		normal_cell_26_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,45),
			fetch              => s_fetch(26,45),
			data_in            => s_data_in(26,45),
			data_out           => s_data_out(26,45),
			out1               => s_out1(26,45),
			out2               => s_out2(26,45),
			lock_lower_row_out => s_locks_lower_out(26,45),
			lock_lower_row_in  => s_locks_lower_in(26,45),
			in1                => s_in1(26,45),
			in2                => s_in2(26,45),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(45)
		);
	s_in1(26,45)            <= s_out1(27,45);
	s_in2(26,45)            <= s_out2(27,46);
	s_locks_lower_in(26,45) <= s_locks_lower_out(27,45);

		normal_cell_26_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,46),
			fetch              => s_fetch(26,46),
			data_in            => s_data_in(26,46),
			data_out           => s_data_out(26,46),
			out1               => s_out1(26,46),
			out2               => s_out2(26,46),
			lock_lower_row_out => s_locks_lower_out(26,46),
			lock_lower_row_in  => s_locks_lower_in(26,46),
			in1                => s_in1(26,46),
			in2                => s_in2(26,46),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(46)
		);
	s_in1(26,46)            <= s_out1(27,46);
	s_in2(26,46)            <= s_out2(27,47);
	s_locks_lower_in(26,46) <= s_locks_lower_out(27,46);

		normal_cell_26_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,47),
			fetch              => s_fetch(26,47),
			data_in            => s_data_in(26,47),
			data_out           => s_data_out(26,47),
			out1               => s_out1(26,47),
			out2               => s_out2(26,47),
			lock_lower_row_out => s_locks_lower_out(26,47),
			lock_lower_row_in  => s_locks_lower_in(26,47),
			in1                => s_in1(26,47),
			in2                => s_in2(26,47),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(47)
		);
	s_in1(26,47)            <= s_out1(27,47);
	s_in2(26,47)            <= s_out2(27,48);
	s_locks_lower_in(26,47) <= s_locks_lower_out(27,47);

		normal_cell_26_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,48),
			fetch              => s_fetch(26,48),
			data_in            => s_data_in(26,48),
			data_out           => s_data_out(26,48),
			out1               => s_out1(26,48),
			out2               => s_out2(26,48),
			lock_lower_row_out => s_locks_lower_out(26,48),
			lock_lower_row_in  => s_locks_lower_in(26,48),
			in1                => s_in1(26,48),
			in2                => s_in2(26,48),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(48)
		);
	s_in1(26,48)            <= s_out1(27,48);
	s_in2(26,48)            <= s_out2(27,49);
	s_locks_lower_in(26,48) <= s_locks_lower_out(27,48);

		normal_cell_26_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,49),
			fetch              => s_fetch(26,49),
			data_in            => s_data_in(26,49),
			data_out           => s_data_out(26,49),
			out1               => s_out1(26,49),
			out2               => s_out2(26,49),
			lock_lower_row_out => s_locks_lower_out(26,49),
			lock_lower_row_in  => s_locks_lower_in(26,49),
			in1                => s_in1(26,49),
			in2                => s_in2(26,49),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(49)
		);
	s_in1(26,49)            <= s_out1(27,49);
	s_in2(26,49)            <= s_out2(27,50);
	s_locks_lower_in(26,49) <= s_locks_lower_out(27,49);

		normal_cell_26_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,50),
			fetch              => s_fetch(26,50),
			data_in            => s_data_in(26,50),
			data_out           => s_data_out(26,50),
			out1               => s_out1(26,50),
			out2               => s_out2(26,50),
			lock_lower_row_out => s_locks_lower_out(26,50),
			lock_lower_row_in  => s_locks_lower_in(26,50),
			in1                => s_in1(26,50),
			in2                => s_in2(26,50),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(50)
		);
	s_in1(26,50)            <= s_out1(27,50);
	s_in2(26,50)            <= s_out2(27,51);
	s_locks_lower_in(26,50) <= s_locks_lower_out(27,50);

		normal_cell_26_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,51),
			fetch              => s_fetch(26,51),
			data_in            => s_data_in(26,51),
			data_out           => s_data_out(26,51),
			out1               => s_out1(26,51),
			out2               => s_out2(26,51),
			lock_lower_row_out => s_locks_lower_out(26,51),
			lock_lower_row_in  => s_locks_lower_in(26,51),
			in1                => s_in1(26,51),
			in2                => s_in2(26,51),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(51)
		);
	s_in1(26,51)            <= s_out1(27,51);
	s_in2(26,51)            <= s_out2(27,52);
	s_locks_lower_in(26,51) <= s_locks_lower_out(27,51);

		normal_cell_26_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,52),
			fetch              => s_fetch(26,52),
			data_in            => s_data_in(26,52),
			data_out           => s_data_out(26,52),
			out1               => s_out1(26,52),
			out2               => s_out2(26,52),
			lock_lower_row_out => s_locks_lower_out(26,52),
			lock_lower_row_in  => s_locks_lower_in(26,52),
			in1                => s_in1(26,52),
			in2                => s_in2(26,52),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(52)
		);
	s_in1(26,52)            <= s_out1(27,52);
	s_in2(26,52)            <= s_out2(27,53);
	s_locks_lower_in(26,52) <= s_locks_lower_out(27,52);

		normal_cell_26_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,53),
			fetch              => s_fetch(26,53),
			data_in            => s_data_in(26,53),
			data_out           => s_data_out(26,53),
			out1               => s_out1(26,53),
			out2               => s_out2(26,53),
			lock_lower_row_out => s_locks_lower_out(26,53),
			lock_lower_row_in  => s_locks_lower_in(26,53),
			in1                => s_in1(26,53),
			in2                => s_in2(26,53),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(53)
		);
	s_in1(26,53)            <= s_out1(27,53);
	s_in2(26,53)            <= s_out2(27,54);
	s_locks_lower_in(26,53) <= s_locks_lower_out(27,53);

		normal_cell_26_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,54),
			fetch              => s_fetch(26,54),
			data_in            => s_data_in(26,54),
			data_out           => s_data_out(26,54),
			out1               => s_out1(26,54),
			out2               => s_out2(26,54),
			lock_lower_row_out => s_locks_lower_out(26,54),
			lock_lower_row_in  => s_locks_lower_in(26,54),
			in1                => s_in1(26,54),
			in2                => s_in2(26,54),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(54)
		);
	s_in1(26,54)            <= s_out1(27,54);
	s_in2(26,54)            <= s_out2(27,55);
	s_locks_lower_in(26,54) <= s_locks_lower_out(27,54);

		normal_cell_26_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,55),
			fetch              => s_fetch(26,55),
			data_in            => s_data_in(26,55),
			data_out           => s_data_out(26,55),
			out1               => s_out1(26,55),
			out2               => s_out2(26,55),
			lock_lower_row_out => s_locks_lower_out(26,55),
			lock_lower_row_in  => s_locks_lower_in(26,55),
			in1                => s_in1(26,55),
			in2                => s_in2(26,55),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(55)
		);
	s_in1(26,55)            <= s_out1(27,55);
	s_in2(26,55)            <= s_out2(27,56);
	s_locks_lower_in(26,55) <= s_locks_lower_out(27,55);

		normal_cell_26_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,56),
			fetch              => s_fetch(26,56),
			data_in            => s_data_in(26,56),
			data_out           => s_data_out(26,56),
			out1               => s_out1(26,56),
			out2               => s_out2(26,56),
			lock_lower_row_out => s_locks_lower_out(26,56),
			lock_lower_row_in  => s_locks_lower_in(26,56),
			in1                => s_in1(26,56),
			in2                => s_in2(26,56),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(56)
		);
	s_in1(26,56)            <= s_out1(27,56);
	s_in2(26,56)            <= s_out2(27,57);
	s_locks_lower_in(26,56) <= s_locks_lower_out(27,56);

		normal_cell_26_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,57),
			fetch              => s_fetch(26,57),
			data_in            => s_data_in(26,57),
			data_out           => s_data_out(26,57),
			out1               => s_out1(26,57),
			out2               => s_out2(26,57),
			lock_lower_row_out => s_locks_lower_out(26,57),
			lock_lower_row_in  => s_locks_lower_in(26,57),
			in1                => s_in1(26,57),
			in2                => s_in2(26,57),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(57)
		);
	s_in1(26,57)            <= s_out1(27,57);
	s_in2(26,57)            <= s_out2(27,58);
	s_locks_lower_in(26,57) <= s_locks_lower_out(27,57);

		normal_cell_26_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,58),
			fetch              => s_fetch(26,58),
			data_in            => s_data_in(26,58),
			data_out           => s_data_out(26,58),
			out1               => s_out1(26,58),
			out2               => s_out2(26,58),
			lock_lower_row_out => s_locks_lower_out(26,58),
			lock_lower_row_in  => s_locks_lower_in(26,58),
			in1                => s_in1(26,58),
			in2                => s_in2(26,58),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(58)
		);
	s_in1(26,58)            <= s_out1(27,58);
	s_in2(26,58)            <= s_out2(27,59);
	s_locks_lower_in(26,58) <= s_locks_lower_out(27,58);

		normal_cell_26_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,59),
			fetch              => s_fetch(26,59),
			data_in            => s_data_in(26,59),
			data_out           => s_data_out(26,59),
			out1               => s_out1(26,59),
			out2               => s_out2(26,59),
			lock_lower_row_out => s_locks_lower_out(26,59),
			lock_lower_row_in  => s_locks_lower_in(26,59),
			in1                => s_in1(26,59),
			in2                => s_in2(26,59),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(59)
		);
	s_in1(26,59)            <= s_out1(27,59);
	s_in2(26,59)            <= s_out2(27,60);
	s_locks_lower_in(26,59) <= s_locks_lower_out(27,59);

		last_col_cell_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(26,60),
			fetch              => s_fetch(26,60),
			data_in            => s_data_in(26,60),
			data_out           => s_data_out(26,60),
			out1               => s_out1(26,60),
			out2               => s_out2(26,60),
			lock_lower_row_out => s_locks_lower_out(26,60),
			lock_lower_row_in  => s_locks_lower_in(26,60),
			in1                => s_in1(26,60),
			in2                => (others => '0'),
			lock_row           => s_locks(26),
			piv_found          => s_piv_found,
			row_data           => s_row_data(26),
			col_data           => s_col_data(60)
		);
	s_in1(26,60)            <= s_out1(27,60);
	s_locks_lower_in(26,60) <= s_locks_lower_out(27,60);

		normal_cell_27_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,1),
			fetch              => s_fetch(27,1),
			data_in            => s_data_in(27,1),
			data_out           => s_data_out(27,1),
			out1               => s_out1(27,1),
			out2               => s_out2(27,1),
			lock_lower_row_out => s_locks_lower_out(27,1),
			lock_lower_row_in  => s_locks_lower_in(27,1),
			in1                => s_in1(27,1),
			in2                => s_in2(27,1),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(1)
		);
	s_in1(27,1)            <= s_out1(28,1);
	s_in2(27,1)            <= s_out2(28,2);
	s_locks_lower_in(27,1) <= s_locks_lower_out(28,1);

		normal_cell_27_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,2),
			fetch              => s_fetch(27,2),
			data_in            => s_data_in(27,2),
			data_out           => s_data_out(27,2),
			out1               => s_out1(27,2),
			out2               => s_out2(27,2),
			lock_lower_row_out => s_locks_lower_out(27,2),
			lock_lower_row_in  => s_locks_lower_in(27,2),
			in1                => s_in1(27,2),
			in2                => s_in2(27,2),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(2)
		);
	s_in1(27,2)            <= s_out1(28,2);
	s_in2(27,2)            <= s_out2(28,3);
	s_locks_lower_in(27,2) <= s_locks_lower_out(28,2);

		normal_cell_27_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,3),
			fetch              => s_fetch(27,3),
			data_in            => s_data_in(27,3),
			data_out           => s_data_out(27,3),
			out1               => s_out1(27,3),
			out2               => s_out2(27,3),
			lock_lower_row_out => s_locks_lower_out(27,3),
			lock_lower_row_in  => s_locks_lower_in(27,3),
			in1                => s_in1(27,3),
			in2                => s_in2(27,3),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(3)
		);
	s_in1(27,3)            <= s_out1(28,3);
	s_in2(27,3)            <= s_out2(28,4);
	s_locks_lower_in(27,3) <= s_locks_lower_out(28,3);

		normal_cell_27_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,4),
			fetch              => s_fetch(27,4),
			data_in            => s_data_in(27,4),
			data_out           => s_data_out(27,4),
			out1               => s_out1(27,4),
			out2               => s_out2(27,4),
			lock_lower_row_out => s_locks_lower_out(27,4),
			lock_lower_row_in  => s_locks_lower_in(27,4),
			in1                => s_in1(27,4),
			in2                => s_in2(27,4),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(4)
		);
	s_in1(27,4)            <= s_out1(28,4);
	s_in2(27,4)            <= s_out2(28,5);
	s_locks_lower_in(27,4) <= s_locks_lower_out(28,4);

		normal_cell_27_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,5),
			fetch              => s_fetch(27,5),
			data_in            => s_data_in(27,5),
			data_out           => s_data_out(27,5),
			out1               => s_out1(27,5),
			out2               => s_out2(27,5),
			lock_lower_row_out => s_locks_lower_out(27,5),
			lock_lower_row_in  => s_locks_lower_in(27,5),
			in1                => s_in1(27,5),
			in2                => s_in2(27,5),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(5)
		);
	s_in1(27,5)            <= s_out1(28,5);
	s_in2(27,5)            <= s_out2(28,6);
	s_locks_lower_in(27,5) <= s_locks_lower_out(28,5);

		normal_cell_27_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,6),
			fetch              => s_fetch(27,6),
			data_in            => s_data_in(27,6),
			data_out           => s_data_out(27,6),
			out1               => s_out1(27,6),
			out2               => s_out2(27,6),
			lock_lower_row_out => s_locks_lower_out(27,6),
			lock_lower_row_in  => s_locks_lower_in(27,6),
			in1                => s_in1(27,6),
			in2                => s_in2(27,6),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(6)
		);
	s_in1(27,6)            <= s_out1(28,6);
	s_in2(27,6)            <= s_out2(28,7);
	s_locks_lower_in(27,6) <= s_locks_lower_out(28,6);

		normal_cell_27_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,7),
			fetch              => s_fetch(27,7),
			data_in            => s_data_in(27,7),
			data_out           => s_data_out(27,7),
			out1               => s_out1(27,7),
			out2               => s_out2(27,7),
			lock_lower_row_out => s_locks_lower_out(27,7),
			lock_lower_row_in  => s_locks_lower_in(27,7),
			in1                => s_in1(27,7),
			in2                => s_in2(27,7),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(7)
		);
	s_in1(27,7)            <= s_out1(28,7);
	s_in2(27,7)            <= s_out2(28,8);
	s_locks_lower_in(27,7) <= s_locks_lower_out(28,7);

		normal_cell_27_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,8),
			fetch              => s_fetch(27,8),
			data_in            => s_data_in(27,8),
			data_out           => s_data_out(27,8),
			out1               => s_out1(27,8),
			out2               => s_out2(27,8),
			lock_lower_row_out => s_locks_lower_out(27,8),
			lock_lower_row_in  => s_locks_lower_in(27,8),
			in1                => s_in1(27,8),
			in2                => s_in2(27,8),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(8)
		);
	s_in1(27,8)            <= s_out1(28,8);
	s_in2(27,8)            <= s_out2(28,9);
	s_locks_lower_in(27,8) <= s_locks_lower_out(28,8);

		normal_cell_27_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,9),
			fetch              => s_fetch(27,9),
			data_in            => s_data_in(27,9),
			data_out           => s_data_out(27,9),
			out1               => s_out1(27,9),
			out2               => s_out2(27,9),
			lock_lower_row_out => s_locks_lower_out(27,9),
			lock_lower_row_in  => s_locks_lower_in(27,9),
			in1                => s_in1(27,9),
			in2                => s_in2(27,9),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(9)
		);
	s_in1(27,9)            <= s_out1(28,9);
	s_in2(27,9)            <= s_out2(28,10);
	s_locks_lower_in(27,9) <= s_locks_lower_out(28,9);

		normal_cell_27_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,10),
			fetch              => s_fetch(27,10),
			data_in            => s_data_in(27,10),
			data_out           => s_data_out(27,10),
			out1               => s_out1(27,10),
			out2               => s_out2(27,10),
			lock_lower_row_out => s_locks_lower_out(27,10),
			lock_lower_row_in  => s_locks_lower_in(27,10),
			in1                => s_in1(27,10),
			in2                => s_in2(27,10),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(10)
		);
	s_in1(27,10)            <= s_out1(28,10);
	s_in2(27,10)            <= s_out2(28,11);
	s_locks_lower_in(27,10) <= s_locks_lower_out(28,10);

		normal_cell_27_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,11),
			fetch              => s_fetch(27,11),
			data_in            => s_data_in(27,11),
			data_out           => s_data_out(27,11),
			out1               => s_out1(27,11),
			out2               => s_out2(27,11),
			lock_lower_row_out => s_locks_lower_out(27,11),
			lock_lower_row_in  => s_locks_lower_in(27,11),
			in1                => s_in1(27,11),
			in2                => s_in2(27,11),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(11)
		);
	s_in1(27,11)            <= s_out1(28,11);
	s_in2(27,11)            <= s_out2(28,12);
	s_locks_lower_in(27,11) <= s_locks_lower_out(28,11);

		normal_cell_27_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,12),
			fetch              => s_fetch(27,12),
			data_in            => s_data_in(27,12),
			data_out           => s_data_out(27,12),
			out1               => s_out1(27,12),
			out2               => s_out2(27,12),
			lock_lower_row_out => s_locks_lower_out(27,12),
			lock_lower_row_in  => s_locks_lower_in(27,12),
			in1                => s_in1(27,12),
			in2                => s_in2(27,12),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(12)
		);
	s_in1(27,12)            <= s_out1(28,12);
	s_in2(27,12)            <= s_out2(28,13);
	s_locks_lower_in(27,12) <= s_locks_lower_out(28,12);

		normal_cell_27_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,13),
			fetch              => s_fetch(27,13),
			data_in            => s_data_in(27,13),
			data_out           => s_data_out(27,13),
			out1               => s_out1(27,13),
			out2               => s_out2(27,13),
			lock_lower_row_out => s_locks_lower_out(27,13),
			lock_lower_row_in  => s_locks_lower_in(27,13),
			in1                => s_in1(27,13),
			in2                => s_in2(27,13),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(13)
		);
	s_in1(27,13)            <= s_out1(28,13);
	s_in2(27,13)            <= s_out2(28,14);
	s_locks_lower_in(27,13) <= s_locks_lower_out(28,13);

		normal_cell_27_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,14),
			fetch              => s_fetch(27,14),
			data_in            => s_data_in(27,14),
			data_out           => s_data_out(27,14),
			out1               => s_out1(27,14),
			out2               => s_out2(27,14),
			lock_lower_row_out => s_locks_lower_out(27,14),
			lock_lower_row_in  => s_locks_lower_in(27,14),
			in1                => s_in1(27,14),
			in2                => s_in2(27,14),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(14)
		);
	s_in1(27,14)            <= s_out1(28,14);
	s_in2(27,14)            <= s_out2(28,15);
	s_locks_lower_in(27,14) <= s_locks_lower_out(28,14);

		normal_cell_27_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,15),
			fetch              => s_fetch(27,15),
			data_in            => s_data_in(27,15),
			data_out           => s_data_out(27,15),
			out1               => s_out1(27,15),
			out2               => s_out2(27,15),
			lock_lower_row_out => s_locks_lower_out(27,15),
			lock_lower_row_in  => s_locks_lower_in(27,15),
			in1                => s_in1(27,15),
			in2                => s_in2(27,15),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(15)
		);
	s_in1(27,15)            <= s_out1(28,15);
	s_in2(27,15)            <= s_out2(28,16);
	s_locks_lower_in(27,15) <= s_locks_lower_out(28,15);

		normal_cell_27_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,16),
			fetch              => s_fetch(27,16),
			data_in            => s_data_in(27,16),
			data_out           => s_data_out(27,16),
			out1               => s_out1(27,16),
			out2               => s_out2(27,16),
			lock_lower_row_out => s_locks_lower_out(27,16),
			lock_lower_row_in  => s_locks_lower_in(27,16),
			in1                => s_in1(27,16),
			in2                => s_in2(27,16),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(16)
		);
	s_in1(27,16)            <= s_out1(28,16);
	s_in2(27,16)            <= s_out2(28,17);
	s_locks_lower_in(27,16) <= s_locks_lower_out(28,16);

		normal_cell_27_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,17),
			fetch              => s_fetch(27,17),
			data_in            => s_data_in(27,17),
			data_out           => s_data_out(27,17),
			out1               => s_out1(27,17),
			out2               => s_out2(27,17),
			lock_lower_row_out => s_locks_lower_out(27,17),
			lock_lower_row_in  => s_locks_lower_in(27,17),
			in1                => s_in1(27,17),
			in2                => s_in2(27,17),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(17)
		);
	s_in1(27,17)            <= s_out1(28,17);
	s_in2(27,17)            <= s_out2(28,18);
	s_locks_lower_in(27,17) <= s_locks_lower_out(28,17);

		normal_cell_27_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,18),
			fetch              => s_fetch(27,18),
			data_in            => s_data_in(27,18),
			data_out           => s_data_out(27,18),
			out1               => s_out1(27,18),
			out2               => s_out2(27,18),
			lock_lower_row_out => s_locks_lower_out(27,18),
			lock_lower_row_in  => s_locks_lower_in(27,18),
			in1                => s_in1(27,18),
			in2                => s_in2(27,18),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(18)
		);
	s_in1(27,18)            <= s_out1(28,18);
	s_in2(27,18)            <= s_out2(28,19);
	s_locks_lower_in(27,18) <= s_locks_lower_out(28,18);

		normal_cell_27_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,19),
			fetch              => s_fetch(27,19),
			data_in            => s_data_in(27,19),
			data_out           => s_data_out(27,19),
			out1               => s_out1(27,19),
			out2               => s_out2(27,19),
			lock_lower_row_out => s_locks_lower_out(27,19),
			lock_lower_row_in  => s_locks_lower_in(27,19),
			in1                => s_in1(27,19),
			in2                => s_in2(27,19),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(19)
		);
	s_in1(27,19)            <= s_out1(28,19);
	s_in2(27,19)            <= s_out2(28,20);
	s_locks_lower_in(27,19) <= s_locks_lower_out(28,19);

		normal_cell_27_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,20),
			fetch              => s_fetch(27,20),
			data_in            => s_data_in(27,20),
			data_out           => s_data_out(27,20),
			out1               => s_out1(27,20),
			out2               => s_out2(27,20),
			lock_lower_row_out => s_locks_lower_out(27,20),
			lock_lower_row_in  => s_locks_lower_in(27,20),
			in1                => s_in1(27,20),
			in2                => s_in2(27,20),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(20)
		);
	s_in1(27,20)            <= s_out1(28,20);
	s_in2(27,20)            <= s_out2(28,21);
	s_locks_lower_in(27,20) <= s_locks_lower_out(28,20);

		normal_cell_27_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,21),
			fetch              => s_fetch(27,21),
			data_in            => s_data_in(27,21),
			data_out           => s_data_out(27,21),
			out1               => s_out1(27,21),
			out2               => s_out2(27,21),
			lock_lower_row_out => s_locks_lower_out(27,21),
			lock_lower_row_in  => s_locks_lower_in(27,21),
			in1                => s_in1(27,21),
			in2                => s_in2(27,21),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(21)
		);
	s_in1(27,21)            <= s_out1(28,21);
	s_in2(27,21)            <= s_out2(28,22);
	s_locks_lower_in(27,21) <= s_locks_lower_out(28,21);

		normal_cell_27_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,22),
			fetch              => s_fetch(27,22),
			data_in            => s_data_in(27,22),
			data_out           => s_data_out(27,22),
			out1               => s_out1(27,22),
			out2               => s_out2(27,22),
			lock_lower_row_out => s_locks_lower_out(27,22),
			lock_lower_row_in  => s_locks_lower_in(27,22),
			in1                => s_in1(27,22),
			in2                => s_in2(27,22),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(22)
		);
	s_in1(27,22)            <= s_out1(28,22);
	s_in2(27,22)            <= s_out2(28,23);
	s_locks_lower_in(27,22) <= s_locks_lower_out(28,22);

		normal_cell_27_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,23),
			fetch              => s_fetch(27,23),
			data_in            => s_data_in(27,23),
			data_out           => s_data_out(27,23),
			out1               => s_out1(27,23),
			out2               => s_out2(27,23),
			lock_lower_row_out => s_locks_lower_out(27,23),
			lock_lower_row_in  => s_locks_lower_in(27,23),
			in1                => s_in1(27,23),
			in2                => s_in2(27,23),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(23)
		);
	s_in1(27,23)            <= s_out1(28,23);
	s_in2(27,23)            <= s_out2(28,24);
	s_locks_lower_in(27,23) <= s_locks_lower_out(28,23);

		normal_cell_27_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,24),
			fetch              => s_fetch(27,24),
			data_in            => s_data_in(27,24),
			data_out           => s_data_out(27,24),
			out1               => s_out1(27,24),
			out2               => s_out2(27,24),
			lock_lower_row_out => s_locks_lower_out(27,24),
			lock_lower_row_in  => s_locks_lower_in(27,24),
			in1                => s_in1(27,24),
			in2                => s_in2(27,24),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(24)
		);
	s_in1(27,24)            <= s_out1(28,24);
	s_in2(27,24)            <= s_out2(28,25);
	s_locks_lower_in(27,24) <= s_locks_lower_out(28,24);

		normal_cell_27_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,25),
			fetch              => s_fetch(27,25),
			data_in            => s_data_in(27,25),
			data_out           => s_data_out(27,25),
			out1               => s_out1(27,25),
			out2               => s_out2(27,25),
			lock_lower_row_out => s_locks_lower_out(27,25),
			lock_lower_row_in  => s_locks_lower_in(27,25),
			in1                => s_in1(27,25),
			in2                => s_in2(27,25),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(25)
		);
	s_in1(27,25)            <= s_out1(28,25);
	s_in2(27,25)            <= s_out2(28,26);
	s_locks_lower_in(27,25) <= s_locks_lower_out(28,25);

		normal_cell_27_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,26),
			fetch              => s_fetch(27,26),
			data_in            => s_data_in(27,26),
			data_out           => s_data_out(27,26),
			out1               => s_out1(27,26),
			out2               => s_out2(27,26),
			lock_lower_row_out => s_locks_lower_out(27,26),
			lock_lower_row_in  => s_locks_lower_in(27,26),
			in1                => s_in1(27,26),
			in2                => s_in2(27,26),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(26)
		);
	s_in1(27,26)            <= s_out1(28,26);
	s_in2(27,26)            <= s_out2(28,27);
	s_locks_lower_in(27,26) <= s_locks_lower_out(28,26);

		normal_cell_27_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,27),
			fetch              => s_fetch(27,27),
			data_in            => s_data_in(27,27),
			data_out           => s_data_out(27,27),
			out1               => s_out1(27,27),
			out2               => s_out2(27,27),
			lock_lower_row_out => s_locks_lower_out(27,27),
			lock_lower_row_in  => s_locks_lower_in(27,27),
			in1                => s_in1(27,27),
			in2                => s_in2(27,27),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(27)
		);
	s_in1(27,27)            <= s_out1(28,27);
	s_in2(27,27)            <= s_out2(28,28);
	s_locks_lower_in(27,27) <= s_locks_lower_out(28,27);

		normal_cell_27_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,28),
			fetch              => s_fetch(27,28),
			data_in            => s_data_in(27,28),
			data_out           => s_data_out(27,28),
			out1               => s_out1(27,28),
			out2               => s_out2(27,28),
			lock_lower_row_out => s_locks_lower_out(27,28),
			lock_lower_row_in  => s_locks_lower_in(27,28),
			in1                => s_in1(27,28),
			in2                => s_in2(27,28),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(28)
		);
	s_in1(27,28)            <= s_out1(28,28);
	s_in2(27,28)            <= s_out2(28,29);
	s_locks_lower_in(27,28) <= s_locks_lower_out(28,28);

		normal_cell_27_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,29),
			fetch              => s_fetch(27,29),
			data_in            => s_data_in(27,29),
			data_out           => s_data_out(27,29),
			out1               => s_out1(27,29),
			out2               => s_out2(27,29),
			lock_lower_row_out => s_locks_lower_out(27,29),
			lock_lower_row_in  => s_locks_lower_in(27,29),
			in1                => s_in1(27,29),
			in2                => s_in2(27,29),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(29)
		);
	s_in1(27,29)            <= s_out1(28,29);
	s_in2(27,29)            <= s_out2(28,30);
	s_locks_lower_in(27,29) <= s_locks_lower_out(28,29);

		normal_cell_27_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,30),
			fetch              => s_fetch(27,30),
			data_in            => s_data_in(27,30),
			data_out           => s_data_out(27,30),
			out1               => s_out1(27,30),
			out2               => s_out2(27,30),
			lock_lower_row_out => s_locks_lower_out(27,30),
			lock_lower_row_in  => s_locks_lower_in(27,30),
			in1                => s_in1(27,30),
			in2                => s_in2(27,30),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(30)
		);
	s_in1(27,30)            <= s_out1(28,30);
	s_in2(27,30)            <= s_out2(28,31);
	s_locks_lower_in(27,30) <= s_locks_lower_out(28,30);

		normal_cell_27_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,31),
			fetch              => s_fetch(27,31),
			data_in            => s_data_in(27,31),
			data_out           => s_data_out(27,31),
			out1               => s_out1(27,31),
			out2               => s_out2(27,31),
			lock_lower_row_out => s_locks_lower_out(27,31),
			lock_lower_row_in  => s_locks_lower_in(27,31),
			in1                => s_in1(27,31),
			in2                => s_in2(27,31),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(31)
		);
	s_in1(27,31)            <= s_out1(28,31);
	s_in2(27,31)            <= s_out2(28,32);
	s_locks_lower_in(27,31) <= s_locks_lower_out(28,31);

		normal_cell_27_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,32),
			fetch              => s_fetch(27,32),
			data_in            => s_data_in(27,32),
			data_out           => s_data_out(27,32),
			out1               => s_out1(27,32),
			out2               => s_out2(27,32),
			lock_lower_row_out => s_locks_lower_out(27,32),
			lock_lower_row_in  => s_locks_lower_in(27,32),
			in1                => s_in1(27,32),
			in2                => s_in2(27,32),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(32)
		);
	s_in1(27,32)            <= s_out1(28,32);
	s_in2(27,32)            <= s_out2(28,33);
	s_locks_lower_in(27,32) <= s_locks_lower_out(28,32);

		normal_cell_27_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,33),
			fetch              => s_fetch(27,33),
			data_in            => s_data_in(27,33),
			data_out           => s_data_out(27,33),
			out1               => s_out1(27,33),
			out2               => s_out2(27,33),
			lock_lower_row_out => s_locks_lower_out(27,33),
			lock_lower_row_in  => s_locks_lower_in(27,33),
			in1                => s_in1(27,33),
			in2                => s_in2(27,33),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(33)
		);
	s_in1(27,33)            <= s_out1(28,33);
	s_in2(27,33)            <= s_out2(28,34);
	s_locks_lower_in(27,33) <= s_locks_lower_out(28,33);

		normal_cell_27_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,34),
			fetch              => s_fetch(27,34),
			data_in            => s_data_in(27,34),
			data_out           => s_data_out(27,34),
			out1               => s_out1(27,34),
			out2               => s_out2(27,34),
			lock_lower_row_out => s_locks_lower_out(27,34),
			lock_lower_row_in  => s_locks_lower_in(27,34),
			in1                => s_in1(27,34),
			in2                => s_in2(27,34),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(34)
		);
	s_in1(27,34)            <= s_out1(28,34);
	s_in2(27,34)            <= s_out2(28,35);
	s_locks_lower_in(27,34) <= s_locks_lower_out(28,34);

		normal_cell_27_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,35),
			fetch              => s_fetch(27,35),
			data_in            => s_data_in(27,35),
			data_out           => s_data_out(27,35),
			out1               => s_out1(27,35),
			out2               => s_out2(27,35),
			lock_lower_row_out => s_locks_lower_out(27,35),
			lock_lower_row_in  => s_locks_lower_in(27,35),
			in1                => s_in1(27,35),
			in2                => s_in2(27,35),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(35)
		);
	s_in1(27,35)            <= s_out1(28,35);
	s_in2(27,35)            <= s_out2(28,36);
	s_locks_lower_in(27,35) <= s_locks_lower_out(28,35);

		normal_cell_27_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,36),
			fetch              => s_fetch(27,36),
			data_in            => s_data_in(27,36),
			data_out           => s_data_out(27,36),
			out1               => s_out1(27,36),
			out2               => s_out2(27,36),
			lock_lower_row_out => s_locks_lower_out(27,36),
			lock_lower_row_in  => s_locks_lower_in(27,36),
			in1                => s_in1(27,36),
			in2                => s_in2(27,36),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(36)
		);
	s_in1(27,36)            <= s_out1(28,36);
	s_in2(27,36)            <= s_out2(28,37);
	s_locks_lower_in(27,36) <= s_locks_lower_out(28,36);

		normal_cell_27_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,37),
			fetch              => s_fetch(27,37),
			data_in            => s_data_in(27,37),
			data_out           => s_data_out(27,37),
			out1               => s_out1(27,37),
			out2               => s_out2(27,37),
			lock_lower_row_out => s_locks_lower_out(27,37),
			lock_lower_row_in  => s_locks_lower_in(27,37),
			in1                => s_in1(27,37),
			in2                => s_in2(27,37),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(37)
		);
	s_in1(27,37)            <= s_out1(28,37);
	s_in2(27,37)            <= s_out2(28,38);
	s_locks_lower_in(27,37) <= s_locks_lower_out(28,37);

		normal_cell_27_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,38),
			fetch              => s_fetch(27,38),
			data_in            => s_data_in(27,38),
			data_out           => s_data_out(27,38),
			out1               => s_out1(27,38),
			out2               => s_out2(27,38),
			lock_lower_row_out => s_locks_lower_out(27,38),
			lock_lower_row_in  => s_locks_lower_in(27,38),
			in1                => s_in1(27,38),
			in2                => s_in2(27,38),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(38)
		);
	s_in1(27,38)            <= s_out1(28,38);
	s_in2(27,38)            <= s_out2(28,39);
	s_locks_lower_in(27,38) <= s_locks_lower_out(28,38);

		normal_cell_27_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,39),
			fetch              => s_fetch(27,39),
			data_in            => s_data_in(27,39),
			data_out           => s_data_out(27,39),
			out1               => s_out1(27,39),
			out2               => s_out2(27,39),
			lock_lower_row_out => s_locks_lower_out(27,39),
			lock_lower_row_in  => s_locks_lower_in(27,39),
			in1                => s_in1(27,39),
			in2                => s_in2(27,39),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(39)
		);
	s_in1(27,39)            <= s_out1(28,39);
	s_in2(27,39)            <= s_out2(28,40);
	s_locks_lower_in(27,39) <= s_locks_lower_out(28,39);

		normal_cell_27_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,40),
			fetch              => s_fetch(27,40),
			data_in            => s_data_in(27,40),
			data_out           => s_data_out(27,40),
			out1               => s_out1(27,40),
			out2               => s_out2(27,40),
			lock_lower_row_out => s_locks_lower_out(27,40),
			lock_lower_row_in  => s_locks_lower_in(27,40),
			in1                => s_in1(27,40),
			in2                => s_in2(27,40),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(40)
		);
	s_in1(27,40)            <= s_out1(28,40);
	s_in2(27,40)            <= s_out2(28,41);
	s_locks_lower_in(27,40) <= s_locks_lower_out(28,40);

		normal_cell_27_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,41),
			fetch              => s_fetch(27,41),
			data_in            => s_data_in(27,41),
			data_out           => s_data_out(27,41),
			out1               => s_out1(27,41),
			out2               => s_out2(27,41),
			lock_lower_row_out => s_locks_lower_out(27,41),
			lock_lower_row_in  => s_locks_lower_in(27,41),
			in1                => s_in1(27,41),
			in2                => s_in2(27,41),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(41)
		);
	s_in1(27,41)            <= s_out1(28,41);
	s_in2(27,41)            <= s_out2(28,42);
	s_locks_lower_in(27,41) <= s_locks_lower_out(28,41);

		normal_cell_27_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,42),
			fetch              => s_fetch(27,42),
			data_in            => s_data_in(27,42),
			data_out           => s_data_out(27,42),
			out1               => s_out1(27,42),
			out2               => s_out2(27,42),
			lock_lower_row_out => s_locks_lower_out(27,42),
			lock_lower_row_in  => s_locks_lower_in(27,42),
			in1                => s_in1(27,42),
			in2                => s_in2(27,42),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(42)
		);
	s_in1(27,42)            <= s_out1(28,42);
	s_in2(27,42)            <= s_out2(28,43);
	s_locks_lower_in(27,42) <= s_locks_lower_out(28,42);

		normal_cell_27_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,43),
			fetch              => s_fetch(27,43),
			data_in            => s_data_in(27,43),
			data_out           => s_data_out(27,43),
			out1               => s_out1(27,43),
			out2               => s_out2(27,43),
			lock_lower_row_out => s_locks_lower_out(27,43),
			lock_lower_row_in  => s_locks_lower_in(27,43),
			in1                => s_in1(27,43),
			in2                => s_in2(27,43),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(43)
		);
	s_in1(27,43)            <= s_out1(28,43);
	s_in2(27,43)            <= s_out2(28,44);
	s_locks_lower_in(27,43) <= s_locks_lower_out(28,43);

		normal_cell_27_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,44),
			fetch              => s_fetch(27,44),
			data_in            => s_data_in(27,44),
			data_out           => s_data_out(27,44),
			out1               => s_out1(27,44),
			out2               => s_out2(27,44),
			lock_lower_row_out => s_locks_lower_out(27,44),
			lock_lower_row_in  => s_locks_lower_in(27,44),
			in1                => s_in1(27,44),
			in2                => s_in2(27,44),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(44)
		);
	s_in1(27,44)            <= s_out1(28,44);
	s_in2(27,44)            <= s_out2(28,45);
	s_locks_lower_in(27,44) <= s_locks_lower_out(28,44);

		normal_cell_27_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,45),
			fetch              => s_fetch(27,45),
			data_in            => s_data_in(27,45),
			data_out           => s_data_out(27,45),
			out1               => s_out1(27,45),
			out2               => s_out2(27,45),
			lock_lower_row_out => s_locks_lower_out(27,45),
			lock_lower_row_in  => s_locks_lower_in(27,45),
			in1                => s_in1(27,45),
			in2                => s_in2(27,45),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(45)
		);
	s_in1(27,45)            <= s_out1(28,45);
	s_in2(27,45)            <= s_out2(28,46);
	s_locks_lower_in(27,45) <= s_locks_lower_out(28,45);

		normal_cell_27_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,46),
			fetch              => s_fetch(27,46),
			data_in            => s_data_in(27,46),
			data_out           => s_data_out(27,46),
			out1               => s_out1(27,46),
			out2               => s_out2(27,46),
			lock_lower_row_out => s_locks_lower_out(27,46),
			lock_lower_row_in  => s_locks_lower_in(27,46),
			in1                => s_in1(27,46),
			in2                => s_in2(27,46),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(46)
		);
	s_in1(27,46)            <= s_out1(28,46);
	s_in2(27,46)            <= s_out2(28,47);
	s_locks_lower_in(27,46) <= s_locks_lower_out(28,46);

		normal_cell_27_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,47),
			fetch              => s_fetch(27,47),
			data_in            => s_data_in(27,47),
			data_out           => s_data_out(27,47),
			out1               => s_out1(27,47),
			out2               => s_out2(27,47),
			lock_lower_row_out => s_locks_lower_out(27,47),
			lock_lower_row_in  => s_locks_lower_in(27,47),
			in1                => s_in1(27,47),
			in2                => s_in2(27,47),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(47)
		);
	s_in1(27,47)            <= s_out1(28,47);
	s_in2(27,47)            <= s_out2(28,48);
	s_locks_lower_in(27,47) <= s_locks_lower_out(28,47);

		normal_cell_27_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,48),
			fetch              => s_fetch(27,48),
			data_in            => s_data_in(27,48),
			data_out           => s_data_out(27,48),
			out1               => s_out1(27,48),
			out2               => s_out2(27,48),
			lock_lower_row_out => s_locks_lower_out(27,48),
			lock_lower_row_in  => s_locks_lower_in(27,48),
			in1                => s_in1(27,48),
			in2                => s_in2(27,48),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(48)
		);
	s_in1(27,48)            <= s_out1(28,48);
	s_in2(27,48)            <= s_out2(28,49);
	s_locks_lower_in(27,48) <= s_locks_lower_out(28,48);

		normal_cell_27_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,49),
			fetch              => s_fetch(27,49),
			data_in            => s_data_in(27,49),
			data_out           => s_data_out(27,49),
			out1               => s_out1(27,49),
			out2               => s_out2(27,49),
			lock_lower_row_out => s_locks_lower_out(27,49),
			lock_lower_row_in  => s_locks_lower_in(27,49),
			in1                => s_in1(27,49),
			in2                => s_in2(27,49),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(49)
		);
	s_in1(27,49)            <= s_out1(28,49);
	s_in2(27,49)            <= s_out2(28,50);
	s_locks_lower_in(27,49) <= s_locks_lower_out(28,49);

		normal_cell_27_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,50),
			fetch              => s_fetch(27,50),
			data_in            => s_data_in(27,50),
			data_out           => s_data_out(27,50),
			out1               => s_out1(27,50),
			out2               => s_out2(27,50),
			lock_lower_row_out => s_locks_lower_out(27,50),
			lock_lower_row_in  => s_locks_lower_in(27,50),
			in1                => s_in1(27,50),
			in2                => s_in2(27,50),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(50)
		);
	s_in1(27,50)            <= s_out1(28,50);
	s_in2(27,50)            <= s_out2(28,51);
	s_locks_lower_in(27,50) <= s_locks_lower_out(28,50);

		normal_cell_27_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,51),
			fetch              => s_fetch(27,51),
			data_in            => s_data_in(27,51),
			data_out           => s_data_out(27,51),
			out1               => s_out1(27,51),
			out2               => s_out2(27,51),
			lock_lower_row_out => s_locks_lower_out(27,51),
			lock_lower_row_in  => s_locks_lower_in(27,51),
			in1                => s_in1(27,51),
			in2                => s_in2(27,51),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(51)
		);
	s_in1(27,51)            <= s_out1(28,51);
	s_in2(27,51)            <= s_out2(28,52);
	s_locks_lower_in(27,51) <= s_locks_lower_out(28,51);

		normal_cell_27_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,52),
			fetch              => s_fetch(27,52),
			data_in            => s_data_in(27,52),
			data_out           => s_data_out(27,52),
			out1               => s_out1(27,52),
			out2               => s_out2(27,52),
			lock_lower_row_out => s_locks_lower_out(27,52),
			lock_lower_row_in  => s_locks_lower_in(27,52),
			in1                => s_in1(27,52),
			in2                => s_in2(27,52),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(52)
		);
	s_in1(27,52)            <= s_out1(28,52);
	s_in2(27,52)            <= s_out2(28,53);
	s_locks_lower_in(27,52) <= s_locks_lower_out(28,52);

		normal_cell_27_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,53),
			fetch              => s_fetch(27,53),
			data_in            => s_data_in(27,53),
			data_out           => s_data_out(27,53),
			out1               => s_out1(27,53),
			out2               => s_out2(27,53),
			lock_lower_row_out => s_locks_lower_out(27,53),
			lock_lower_row_in  => s_locks_lower_in(27,53),
			in1                => s_in1(27,53),
			in2                => s_in2(27,53),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(53)
		);
	s_in1(27,53)            <= s_out1(28,53);
	s_in2(27,53)            <= s_out2(28,54);
	s_locks_lower_in(27,53) <= s_locks_lower_out(28,53);

		normal_cell_27_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,54),
			fetch              => s_fetch(27,54),
			data_in            => s_data_in(27,54),
			data_out           => s_data_out(27,54),
			out1               => s_out1(27,54),
			out2               => s_out2(27,54),
			lock_lower_row_out => s_locks_lower_out(27,54),
			lock_lower_row_in  => s_locks_lower_in(27,54),
			in1                => s_in1(27,54),
			in2                => s_in2(27,54),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(54)
		);
	s_in1(27,54)            <= s_out1(28,54);
	s_in2(27,54)            <= s_out2(28,55);
	s_locks_lower_in(27,54) <= s_locks_lower_out(28,54);

		normal_cell_27_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,55),
			fetch              => s_fetch(27,55),
			data_in            => s_data_in(27,55),
			data_out           => s_data_out(27,55),
			out1               => s_out1(27,55),
			out2               => s_out2(27,55),
			lock_lower_row_out => s_locks_lower_out(27,55),
			lock_lower_row_in  => s_locks_lower_in(27,55),
			in1                => s_in1(27,55),
			in2                => s_in2(27,55),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(55)
		);
	s_in1(27,55)            <= s_out1(28,55);
	s_in2(27,55)            <= s_out2(28,56);
	s_locks_lower_in(27,55) <= s_locks_lower_out(28,55);

		normal_cell_27_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,56),
			fetch              => s_fetch(27,56),
			data_in            => s_data_in(27,56),
			data_out           => s_data_out(27,56),
			out1               => s_out1(27,56),
			out2               => s_out2(27,56),
			lock_lower_row_out => s_locks_lower_out(27,56),
			lock_lower_row_in  => s_locks_lower_in(27,56),
			in1                => s_in1(27,56),
			in2                => s_in2(27,56),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(56)
		);
	s_in1(27,56)            <= s_out1(28,56);
	s_in2(27,56)            <= s_out2(28,57);
	s_locks_lower_in(27,56) <= s_locks_lower_out(28,56);

		normal_cell_27_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,57),
			fetch              => s_fetch(27,57),
			data_in            => s_data_in(27,57),
			data_out           => s_data_out(27,57),
			out1               => s_out1(27,57),
			out2               => s_out2(27,57),
			lock_lower_row_out => s_locks_lower_out(27,57),
			lock_lower_row_in  => s_locks_lower_in(27,57),
			in1                => s_in1(27,57),
			in2                => s_in2(27,57),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(57)
		);
	s_in1(27,57)            <= s_out1(28,57);
	s_in2(27,57)            <= s_out2(28,58);
	s_locks_lower_in(27,57) <= s_locks_lower_out(28,57);

		normal_cell_27_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,58),
			fetch              => s_fetch(27,58),
			data_in            => s_data_in(27,58),
			data_out           => s_data_out(27,58),
			out1               => s_out1(27,58),
			out2               => s_out2(27,58),
			lock_lower_row_out => s_locks_lower_out(27,58),
			lock_lower_row_in  => s_locks_lower_in(27,58),
			in1                => s_in1(27,58),
			in2                => s_in2(27,58),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(58)
		);
	s_in1(27,58)            <= s_out1(28,58);
	s_in2(27,58)            <= s_out2(28,59);
	s_locks_lower_in(27,58) <= s_locks_lower_out(28,58);

		normal_cell_27_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,59),
			fetch              => s_fetch(27,59),
			data_in            => s_data_in(27,59),
			data_out           => s_data_out(27,59),
			out1               => s_out1(27,59),
			out2               => s_out2(27,59),
			lock_lower_row_out => s_locks_lower_out(27,59),
			lock_lower_row_in  => s_locks_lower_in(27,59),
			in1                => s_in1(27,59),
			in2                => s_in2(27,59),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(59)
		);
	s_in1(27,59)            <= s_out1(28,59);
	s_in2(27,59)            <= s_out2(28,60);
	s_locks_lower_in(27,59) <= s_locks_lower_out(28,59);

		last_col_cell_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(27,60),
			fetch              => s_fetch(27,60),
			data_in            => s_data_in(27,60),
			data_out           => s_data_out(27,60),
			out1               => s_out1(27,60),
			out2               => s_out2(27,60),
			lock_lower_row_out => s_locks_lower_out(27,60),
			lock_lower_row_in  => s_locks_lower_in(27,60),
			in1                => s_in1(27,60),
			in2                => (others => '0'),
			lock_row           => s_locks(27),
			piv_found          => s_piv_found,
			row_data           => s_row_data(27),
			col_data           => s_col_data(60)
		);
	s_in1(27,60)            <= s_out1(28,60);
	s_locks_lower_in(27,60) <= s_locks_lower_out(28,60);

		normal_cell_28_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,1),
			fetch              => s_fetch(28,1),
			data_in            => s_data_in(28,1),
			data_out           => s_data_out(28,1),
			out1               => s_out1(28,1),
			out2               => s_out2(28,1),
			lock_lower_row_out => s_locks_lower_out(28,1),
			lock_lower_row_in  => s_locks_lower_in(28,1),
			in1                => s_in1(28,1),
			in2                => s_in2(28,1),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(1)
		);
	s_in1(28,1)            <= s_out1(29,1);
	s_in2(28,1)            <= s_out2(29,2);
	s_locks_lower_in(28,1) <= s_locks_lower_out(29,1);

		normal_cell_28_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,2),
			fetch              => s_fetch(28,2),
			data_in            => s_data_in(28,2),
			data_out           => s_data_out(28,2),
			out1               => s_out1(28,2),
			out2               => s_out2(28,2),
			lock_lower_row_out => s_locks_lower_out(28,2),
			lock_lower_row_in  => s_locks_lower_in(28,2),
			in1                => s_in1(28,2),
			in2                => s_in2(28,2),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(2)
		);
	s_in1(28,2)            <= s_out1(29,2);
	s_in2(28,2)            <= s_out2(29,3);
	s_locks_lower_in(28,2) <= s_locks_lower_out(29,2);

		normal_cell_28_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,3),
			fetch              => s_fetch(28,3),
			data_in            => s_data_in(28,3),
			data_out           => s_data_out(28,3),
			out1               => s_out1(28,3),
			out2               => s_out2(28,3),
			lock_lower_row_out => s_locks_lower_out(28,3),
			lock_lower_row_in  => s_locks_lower_in(28,3),
			in1                => s_in1(28,3),
			in2                => s_in2(28,3),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(3)
		);
	s_in1(28,3)            <= s_out1(29,3);
	s_in2(28,3)            <= s_out2(29,4);
	s_locks_lower_in(28,3) <= s_locks_lower_out(29,3);

		normal_cell_28_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,4),
			fetch              => s_fetch(28,4),
			data_in            => s_data_in(28,4),
			data_out           => s_data_out(28,4),
			out1               => s_out1(28,4),
			out2               => s_out2(28,4),
			lock_lower_row_out => s_locks_lower_out(28,4),
			lock_lower_row_in  => s_locks_lower_in(28,4),
			in1                => s_in1(28,4),
			in2                => s_in2(28,4),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(4)
		);
	s_in1(28,4)            <= s_out1(29,4);
	s_in2(28,4)            <= s_out2(29,5);
	s_locks_lower_in(28,4) <= s_locks_lower_out(29,4);

		normal_cell_28_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,5),
			fetch              => s_fetch(28,5),
			data_in            => s_data_in(28,5),
			data_out           => s_data_out(28,5),
			out1               => s_out1(28,5),
			out2               => s_out2(28,5),
			lock_lower_row_out => s_locks_lower_out(28,5),
			lock_lower_row_in  => s_locks_lower_in(28,5),
			in1                => s_in1(28,5),
			in2                => s_in2(28,5),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(5)
		);
	s_in1(28,5)            <= s_out1(29,5);
	s_in2(28,5)            <= s_out2(29,6);
	s_locks_lower_in(28,5) <= s_locks_lower_out(29,5);

		normal_cell_28_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,6),
			fetch              => s_fetch(28,6),
			data_in            => s_data_in(28,6),
			data_out           => s_data_out(28,6),
			out1               => s_out1(28,6),
			out2               => s_out2(28,6),
			lock_lower_row_out => s_locks_lower_out(28,6),
			lock_lower_row_in  => s_locks_lower_in(28,6),
			in1                => s_in1(28,6),
			in2                => s_in2(28,6),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(6)
		);
	s_in1(28,6)            <= s_out1(29,6);
	s_in2(28,6)            <= s_out2(29,7);
	s_locks_lower_in(28,6) <= s_locks_lower_out(29,6);

		normal_cell_28_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,7),
			fetch              => s_fetch(28,7),
			data_in            => s_data_in(28,7),
			data_out           => s_data_out(28,7),
			out1               => s_out1(28,7),
			out2               => s_out2(28,7),
			lock_lower_row_out => s_locks_lower_out(28,7),
			lock_lower_row_in  => s_locks_lower_in(28,7),
			in1                => s_in1(28,7),
			in2                => s_in2(28,7),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(7)
		);
	s_in1(28,7)            <= s_out1(29,7);
	s_in2(28,7)            <= s_out2(29,8);
	s_locks_lower_in(28,7) <= s_locks_lower_out(29,7);

		normal_cell_28_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,8),
			fetch              => s_fetch(28,8),
			data_in            => s_data_in(28,8),
			data_out           => s_data_out(28,8),
			out1               => s_out1(28,8),
			out2               => s_out2(28,8),
			lock_lower_row_out => s_locks_lower_out(28,8),
			lock_lower_row_in  => s_locks_lower_in(28,8),
			in1                => s_in1(28,8),
			in2                => s_in2(28,8),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(8)
		);
	s_in1(28,8)            <= s_out1(29,8);
	s_in2(28,8)            <= s_out2(29,9);
	s_locks_lower_in(28,8) <= s_locks_lower_out(29,8);

		normal_cell_28_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,9),
			fetch              => s_fetch(28,9),
			data_in            => s_data_in(28,9),
			data_out           => s_data_out(28,9),
			out1               => s_out1(28,9),
			out2               => s_out2(28,9),
			lock_lower_row_out => s_locks_lower_out(28,9),
			lock_lower_row_in  => s_locks_lower_in(28,9),
			in1                => s_in1(28,9),
			in2                => s_in2(28,9),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(9)
		);
	s_in1(28,9)            <= s_out1(29,9);
	s_in2(28,9)            <= s_out2(29,10);
	s_locks_lower_in(28,9) <= s_locks_lower_out(29,9);

		normal_cell_28_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,10),
			fetch              => s_fetch(28,10),
			data_in            => s_data_in(28,10),
			data_out           => s_data_out(28,10),
			out1               => s_out1(28,10),
			out2               => s_out2(28,10),
			lock_lower_row_out => s_locks_lower_out(28,10),
			lock_lower_row_in  => s_locks_lower_in(28,10),
			in1                => s_in1(28,10),
			in2                => s_in2(28,10),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(10)
		);
	s_in1(28,10)            <= s_out1(29,10);
	s_in2(28,10)            <= s_out2(29,11);
	s_locks_lower_in(28,10) <= s_locks_lower_out(29,10);

		normal_cell_28_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,11),
			fetch              => s_fetch(28,11),
			data_in            => s_data_in(28,11),
			data_out           => s_data_out(28,11),
			out1               => s_out1(28,11),
			out2               => s_out2(28,11),
			lock_lower_row_out => s_locks_lower_out(28,11),
			lock_lower_row_in  => s_locks_lower_in(28,11),
			in1                => s_in1(28,11),
			in2                => s_in2(28,11),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(11)
		);
	s_in1(28,11)            <= s_out1(29,11);
	s_in2(28,11)            <= s_out2(29,12);
	s_locks_lower_in(28,11) <= s_locks_lower_out(29,11);

		normal_cell_28_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,12),
			fetch              => s_fetch(28,12),
			data_in            => s_data_in(28,12),
			data_out           => s_data_out(28,12),
			out1               => s_out1(28,12),
			out2               => s_out2(28,12),
			lock_lower_row_out => s_locks_lower_out(28,12),
			lock_lower_row_in  => s_locks_lower_in(28,12),
			in1                => s_in1(28,12),
			in2                => s_in2(28,12),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(12)
		);
	s_in1(28,12)            <= s_out1(29,12);
	s_in2(28,12)            <= s_out2(29,13);
	s_locks_lower_in(28,12) <= s_locks_lower_out(29,12);

		normal_cell_28_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,13),
			fetch              => s_fetch(28,13),
			data_in            => s_data_in(28,13),
			data_out           => s_data_out(28,13),
			out1               => s_out1(28,13),
			out2               => s_out2(28,13),
			lock_lower_row_out => s_locks_lower_out(28,13),
			lock_lower_row_in  => s_locks_lower_in(28,13),
			in1                => s_in1(28,13),
			in2                => s_in2(28,13),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(13)
		);
	s_in1(28,13)            <= s_out1(29,13);
	s_in2(28,13)            <= s_out2(29,14);
	s_locks_lower_in(28,13) <= s_locks_lower_out(29,13);

		normal_cell_28_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,14),
			fetch              => s_fetch(28,14),
			data_in            => s_data_in(28,14),
			data_out           => s_data_out(28,14),
			out1               => s_out1(28,14),
			out2               => s_out2(28,14),
			lock_lower_row_out => s_locks_lower_out(28,14),
			lock_lower_row_in  => s_locks_lower_in(28,14),
			in1                => s_in1(28,14),
			in2                => s_in2(28,14),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(14)
		);
	s_in1(28,14)            <= s_out1(29,14);
	s_in2(28,14)            <= s_out2(29,15);
	s_locks_lower_in(28,14) <= s_locks_lower_out(29,14);

		normal_cell_28_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,15),
			fetch              => s_fetch(28,15),
			data_in            => s_data_in(28,15),
			data_out           => s_data_out(28,15),
			out1               => s_out1(28,15),
			out2               => s_out2(28,15),
			lock_lower_row_out => s_locks_lower_out(28,15),
			lock_lower_row_in  => s_locks_lower_in(28,15),
			in1                => s_in1(28,15),
			in2                => s_in2(28,15),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(15)
		);
	s_in1(28,15)            <= s_out1(29,15);
	s_in2(28,15)            <= s_out2(29,16);
	s_locks_lower_in(28,15) <= s_locks_lower_out(29,15);

		normal_cell_28_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,16),
			fetch              => s_fetch(28,16),
			data_in            => s_data_in(28,16),
			data_out           => s_data_out(28,16),
			out1               => s_out1(28,16),
			out2               => s_out2(28,16),
			lock_lower_row_out => s_locks_lower_out(28,16),
			lock_lower_row_in  => s_locks_lower_in(28,16),
			in1                => s_in1(28,16),
			in2                => s_in2(28,16),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(16)
		);
	s_in1(28,16)            <= s_out1(29,16);
	s_in2(28,16)            <= s_out2(29,17);
	s_locks_lower_in(28,16) <= s_locks_lower_out(29,16);

		normal_cell_28_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,17),
			fetch              => s_fetch(28,17),
			data_in            => s_data_in(28,17),
			data_out           => s_data_out(28,17),
			out1               => s_out1(28,17),
			out2               => s_out2(28,17),
			lock_lower_row_out => s_locks_lower_out(28,17),
			lock_lower_row_in  => s_locks_lower_in(28,17),
			in1                => s_in1(28,17),
			in2                => s_in2(28,17),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(17)
		);
	s_in1(28,17)            <= s_out1(29,17);
	s_in2(28,17)            <= s_out2(29,18);
	s_locks_lower_in(28,17) <= s_locks_lower_out(29,17);

		normal_cell_28_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,18),
			fetch              => s_fetch(28,18),
			data_in            => s_data_in(28,18),
			data_out           => s_data_out(28,18),
			out1               => s_out1(28,18),
			out2               => s_out2(28,18),
			lock_lower_row_out => s_locks_lower_out(28,18),
			lock_lower_row_in  => s_locks_lower_in(28,18),
			in1                => s_in1(28,18),
			in2                => s_in2(28,18),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(18)
		);
	s_in1(28,18)            <= s_out1(29,18);
	s_in2(28,18)            <= s_out2(29,19);
	s_locks_lower_in(28,18) <= s_locks_lower_out(29,18);

		normal_cell_28_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,19),
			fetch              => s_fetch(28,19),
			data_in            => s_data_in(28,19),
			data_out           => s_data_out(28,19),
			out1               => s_out1(28,19),
			out2               => s_out2(28,19),
			lock_lower_row_out => s_locks_lower_out(28,19),
			lock_lower_row_in  => s_locks_lower_in(28,19),
			in1                => s_in1(28,19),
			in2                => s_in2(28,19),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(19)
		);
	s_in1(28,19)            <= s_out1(29,19);
	s_in2(28,19)            <= s_out2(29,20);
	s_locks_lower_in(28,19) <= s_locks_lower_out(29,19);

		normal_cell_28_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,20),
			fetch              => s_fetch(28,20),
			data_in            => s_data_in(28,20),
			data_out           => s_data_out(28,20),
			out1               => s_out1(28,20),
			out2               => s_out2(28,20),
			lock_lower_row_out => s_locks_lower_out(28,20),
			lock_lower_row_in  => s_locks_lower_in(28,20),
			in1                => s_in1(28,20),
			in2                => s_in2(28,20),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(20)
		);
	s_in1(28,20)            <= s_out1(29,20);
	s_in2(28,20)            <= s_out2(29,21);
	s_locks_lower_in(28,20) <= s_locks_lower_out(29,20);

		normal_cell_28_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,21),
			fetch              => s_fetch(28,21),
			data_in            => s_data_in(28,21),
			data_out           => s_data_out(28,21),
			out1               => s_out1(28,21),
			out2               => s_out2(28,21),
			lock_lower_row_out => s_locks_lower_out(28,21),
			lock_lower_row_in  => s_locks_lower_in(28,21),
			in1                => s_in1(28,21),
			in2                => s_in2(28,21),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(21)
		);
	s_in1(28,21)            <= s_out1(29,21);
	s_in2(28,21)            <= s_out2(29,22);
	s_locks_lower_in(28,21) <= s_locks_lower_out(29,21);

		normal_cell_28_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,22),
			fetch              => s_fetch(28,22),
			data_in            => s_data_in(28,22),
			data_out           => s_data_out(28,22),
			out1               => s_out1(28,22),
			out2               => s_out2(28,22),
			lock_lower_row_out => s_locks_lower_out(28,22),
			lock_lower_row_in  => s_locks_lower_in(28,22),
			in1                => s_in1(28,22),
			in2                => s_in2(28,22),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(22)
		);
	s_in1(28,22)            <= s_out1(29,22);
	s_in2(28,22)            <= s_out2(29,23);
	s_locks_lower_in(28,22) <= s_locks_lower_out(29,22);

		normal_cell_28_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,23),
			fetch              => s_fetch(28,23),
			data_in            => s_data_in(28,23),
			data_out           => s_data_out(28,23),
			out1               => s_out1(28,23),
			out2               => s_out2(28,23),
			lock_lower_row_out => s_locks_lower_out(28,23),
			lock_lower_row_in  => s_locks_lower_in(28,23),
			in1                => s_in1(28,23),
			in2                => s_in2(28,23),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(23)
		);
	s_in1(28,23)            <= s_out1(29,23);
	s_in2(28,23)            <= s_out2(29,24);
	s_locks_lower_in(28,23) <= s_locks_lower_out(29,23);

		normal_cell_28_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,24),
			fetch              => s_fetch(28,24),
			data_in            => s_data_in(28,24),
			data_out           => s_data_out(28,24),
			out1               => s_out1(28,24),
			out2               => s_out2(28,24),
			lock_lower_row_out => s_locks_lower_out(28,24),
			lock_lower_row_in  => s_locks_lower_in(28,24),
			in1                => s_in1(28,24),
			in2                => s_in2(28,24),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(24)
		);
	s_in1(28,24)            <= s_out1(29,24);
	s_in2(28,24)            <= s_out2(29,25);
	s_locks_lower_in(28,24) <= s_locks_lower_out(29,24);

		normal_cell_28_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,25),
			fetch              => s_fetch(28,25),
			data_in            => s_data_in(28,25),
			data_out           => s_data_out(28,25),
			out1               => s_out1(28,25),
			out2               => s_out2(28,25),
			lock_lower_row_out => s_locks_lower_out(28,25),
			lock_lower_row_in  => s_locks_lower_in(28,25),
			in1                => s_in1(28,25),
			in2                => s_in2(28,25),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(25)
		);
	s_in1(28,25)            <= s_out1(29,25);
	s_in2(28,25)            <= s_out2(29,26);
	s_locks_lower_in(28,25) <= s_locks_lower_out(29,25);

		normal_cell_28_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,26),
			fetch              => s_fetch(28,26),
			data_in            => s_data_in(28,26),
			data_out           => s_data_out(28,26),
			out1               => s_out1(28,26),
			out2               => s_out2(28,26),
			lock_lower_row_out => s_locks_lower_out(28,26),
			lock_lower_row_in  => s_locks_lower_in(28,26),
			in1                => s_in1(28,26),
			in2                => s_in2(28,26),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(26)
		);
	s_in1(28,26)            <= s_out1(29,26);
	s_in2(28,26)            <= s_out2(29,27);
	s_locks_lower_in(28,26) <= s_locks_lower_out(29,26);

		normal_cell_28_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,27),
			fetch              => s_fetch(28,27),
			data_in            => s_data_in(28,27),
			data_out           => s_data_out(28,27),
			out1               => s_out1(28,27),
			out2               => s_out2(28,27),
			lock_lower_row_out => s_locks_lower_out(28,27),
			lock_lower_row_in  => s_locks_lower_in(28,27),
			in1                => s_in1(28,27),
			in2                => s_in2(28,27),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(27)
		);
	s_in1(28,27)            <= s_out1(29,27);
	s_in2(28,27)            <= s_out2(29,28);
	s_locks_lower_in(28,27) <= s_locks_lower_out(29,27);

		normal_cell_28_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,28),
			fetch              => s_fetch(28,28),
			data_in            => s_data_in(28,28),
			data_out           => s_data_out(28,28),
			out1               => s_out1(28,28),
			out2               => s_out2(28,28),
			lock_lower_row_out => s_locks_lower_out(28,28),
			lock_lower_row_in  => s_locks_lower_in(28,28),
			in1                => s_in1(28,28),
			in2                => s_in2(28,28),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(28)
		);
	s_in1(28,28)            <= s_out1(29,28);
	s_in2(28,28)            <= s_out2(29,29);
	s_locks_lower_in(28,28) <= s_locks_lower_out(29,28);

		normal_cell_28_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,29),
			fetch              => s_fetch(28,29),
			data_in            => s_data_in(28,29),
			data_out           => s_data_out(28,29),
			out1               => s_out1(28,29),
			out2               => s_out2(28,29),
			lock_lower_row_out => s_locks_lower_out(28,29),
			lock_lower_row_in  => s_locks_lower_in(28,29),
			in1                => s_in1(28,29),
			in2                => s_in2(28,29),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(29)
		);
	s_in1(28,29)            <= s_out1(29,29);
	s_in2(28,29)            <= s_out2(29,30);
	s_locks_lower_in(28,29) <= s_locks_lower_out(29,29);

		normal_cell_28_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,30),
			fetch              => s_fetch(28,30),
			data_in            => s_data_in(28,30),
			data_out           => s_data_out(28,30),
			out1               => s_out1(28,30),
			out2               => s_out2(28,30),
			lock_lower_row_out => s_locks_lower_out(28,30),
			lock_lower_row_in  => s_locks_lower_in(28,30),
			in1                => s_in1(28,30),
			in2                => s_in2(28,30),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(30)
		);
	s_in1(28,30)            <= s_out1(29,30);
	s_in2(28,30)            <= s_out2(29,31);
	s_locks_lower_in(28,30) <= s_locks_lower_out(29,30);

		normal_cell_28_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,31),
			fetch              => s_fetch(28,31),
			data_in            => s_data_in(28,31),
			data_out           => s_data_out(28,31),
			out1               => s_out1(28,31),
			out2               => s_out2(28,31),
			lock_lower_row_out => s_locks_lower_out(28,31),
			lock_lower_row_in  => s_locks_lower_in(28,31),
			in1                => s_in1(28,31),
			in2                => s_in2(28,31),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(31)
		);
	s_in1(28,31)            <= s_out1(29,31);
	s_in2(28,31)            <= s_out2(29,32);
	s_locks_lower_in(28,31) <= s_locks_lower_out(29,31);

		normal_cell_28_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,32),
			fetch              => s_fetch(28,32),
			data_in            => s_data_in(28,32),
			data_out           => s_data_out(28,32),
			out1               => s_out1(28,32),
			out2               => s_out2(28,32),
			lock_lower_row_out => s_locks_lower_out(28,32),
			lock_lower_row_in  => s_locks_lower_in(28,32),
			in1                => s_in1(28,32),
			in2                => s_in2(28,32),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(32)
		);
	s_in1(28,32)            <= s_out1(29,32);
	s_in2(28,32)            <= s_out2(29,33);
	s_locks_lower_in(28,32) <= s_locks_lower_out(29,32);

		normal_cell_28_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,33),
			fetch              => s_fetch(28,33),
			data_in            => s_data_in(28,33),
			data_out           => s_data_out(28,33),
			out1               => s_out1(28,33),
			out2               => s_out2(28,33),
			lock_lower_row_out => s_locks_lower_out(28,33),
			lock_lower_row_in  => s_locks_lower_in(28,33),
			in1                => s_in1(28,33),
			in2                => s_in2(28,33),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(33)
		);
	s_in1(28,33)            <= s_out1(29,33);
	s_in2(28,33)            <= s_out2(29,34);
	s_locks_lower_in(28,33) <= s_locks_lower_out(29,33);

		normal_cell_28_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,34),
			fetch              => s_fetch(28,34),
			data_in            => s_data_in(28,34),
			data_out           => s_data_out(28,34),
			out1               => s_out1(28,34),
			out2               => s_out2(28,34),
			lock_lower_row_out => s_locks_lower_out(28,34),
			lock_lower_row_in  => s_locks_lower_in(28,34),
			in1                => s_in1(28,34),
			in2                => s_in2(28,34),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(34)
		);
	s_in1(28,34)            <= s_out1(29,34);
	s_in2(28,34)            <= s_out2(29,35);
	s_locks_lower_in(28,34) <= s_locks_lower_out(29,34);

		normal_cell_28_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,35),
			fetch              => s_fetch(28,35),
			data_in            => s_data_in(28,35),
			data_out           => s_data_out(28,35),
			out1               => s_out1(28,35),
			out2               => s_out2(28,35),
			lock_lower_row_out => s_locks_lower_out(28,35),
			lock_lower_row_in  => s_locks_lower_in(28,35),
			in1                => s_in1(28,35),
			in2                => s_in2(28,35),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(35)
		);
	s_in1(28,35)            <= s_out1(29,35);
	s_in2(28,35)            <= s_out2(29,36);
	s_locks_lower_in(28,35) <= s_locks_lower_out(29,35);

		normal_cell_28_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,36),
			fetch              => s_fetch(28,36),
			data_in            => s_data_in(28,36),
			data_out           => s_data_out(28,36),
			out1               => s_out1(28,36),
			out2               => s_out2(28,36),
			lock_lower_row_out => s_locks_lower_out(28,36),
			lock_lower_row_in  => s_locks_lower_in(28,36),
			in1                => s_in1(28,36),
			in2                => s_in2(28,36),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(36)
		);
	s_in1(28,36)            <= s_out1(29,36);
	s_in2(28,36)            <= s_out2(29,37);
	s_locks_lower_in(28,36) <= s_locks_lower_out(29,36);

		normal_cell_28_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,37),
			fetch              => s_fetch(28,37),
			data_in            => s_data_in(28,37),
			data_out           => s_data_out(28,37),
			out1               => s_out1(28,37),
			out2               => s_out2(28,37),
			lock_lower_row_out => s_locks_lower_out(28,37),
			lock_lower_row_in  => s_locks_lower_in(28,37),
			in1                => s_in1(28,37),
			in2                => s_in2(28,37),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(37)
		);
	s_in1(28,37)            <= s_out1(29,37);
	s_in2(28,37)            <= s_out2(29,38);
	s_locks_lower_in(28,37) <= s_locks_lower_out(29,37);

		normal_cell_28_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,38),
			fetch              => s_fetch(28,38),
			data_in            => s_data_in(28,38),
			data_out           => s_data_out(28,38),
			out1               => s_out1(28,38),
			out2               => s_out2(28,38),
			lock_lower_row_out => s_locks_lower_out(28,38),
			lock_lower_row_in  => s_locks_lower_in(28,38),
			in1                => s_in1(28,38),
			in2                => s_in2(28,38),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(38)
		);
	s_in1(28,38)            <= s_out1(29,38);
	s_in2(28,38)            <= s_out2(29,39);
	s_locks_lower_in(28,38) <= s_locks_lower_out(29,38);

		normal_cell_28_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,39),
			fetch              => s_fetch(28,39),
			data_in            => s_data_in(28,39),
			data_out           => s_data_out(28,39),
			out1               => s_out1(28,39),
			out2               => s_out2(28,39),
			lock_lower_row_out => s_locks_lower_out(28,39),
			lock_lower_row_in  => s_locks_lower_in(28,39),
			in1                => s_in1(28,39),
			in2                => s_in2(28,39),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(39)
		);
	s_in1(28,39)            <= s_out1(29,39);
	s_in2(28,39)            <= s_out2(29,40);
	s_locks_lower_in(28,39) <= s_locks_lower_out(29,39);

		normal_cell_28_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,40),
			fetch              => s_fetch(28,40),
			data_in            => s_data_in(28,40),
			data_out           => s_data_out(28,40),
			out1               => s_out1(28,40),
			out2               => s_out2(28,40),
			lock_lower_row_out => s_locks_lower_out(28,40),
			lock_lower_row_in  => s_locks_lower_in(28,40),
			in1                => s_in1(28,40),
			in2                => s_in2(28,40),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(40)
		);
	s_in1(28,40)            <= s_out1(29,40);
	s_in2(28,40)            <= s_out2(29,41);
	s_locks_lower_in(28,40) <= s_locks_lower_out(29,40);

		normal_cell_28_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,41),
			fetch              => s_fetch(28,41),
			data_in            => s_data_in(28,41),
			data_out           => s_data_out(28,41),
			out1               => s_out1(28,41),
			out2               => s_out2(28,41),
			lock_lower_row_out => s_locks_lower_out(28,41),
			lock_lower_row_in  => s_locks_lower_in(28,41),
			in1                => s_in1(28,41),
			in2                => s_in2(28,41),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(41)
		);
	s_in1(28,41)            <= s_out1(29,41);
	s_in2(28,41)            <= s_out2(29,42);
	s_locks_lower_in(28,41) <= s_locks_lower_out(29,41);

		normal_cell_28_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,42),
			fetch              => s_fetch(28,42),
			data_in            => s_data_in(28,42),
			data_out           => s_data_out(28,42),
			out1               => s_out1(28,42),
			out2               => s_out2(28,42),
			lock_lower_row_out => s_locks_lower_out(28,42),
			lock_lower_row_in  => s_locks_lower_in(28,42),
			in1                => s_in1(28,42),
			in2                => s_in2(28,42),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(42)
		);
	s_in1(28,42)            <= s_out1(29,42);
	s_in2(28,42)            <= s_out2(29,43);
	s_locks_lower_in(28,42) <= s_locks_lower_out(29,42);

		normal_cell_28_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,43),
			fetch              => s_fetch(28,43),
			data_in            => s_data_in(28,43),
			data_out           => s_data_out(28,43),
			out1               => s_out1(28,43),
			out2               => s_out2(28,43),
			lock_lower_row_out => s_locks_lower_out(28,43),
			lock_lower_row_in  => s_locks_lower_in(28,43),
			in1                => s_in1(28,43),
			in2                => s_in2(28,43),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(43)
		);
	s_in1(28,43)            <= s_out1(29,43);
	s_in2(28,43)            <= s_out2(29,44);
	s_locks_lower_in(28,43) <= s_locks_lower_out(29,43);

		normal_cell_28_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,44),
			fetch              => s_fetch(28,44),
			data_in            => s_data_in(28,44),
			data_out           => s_data_out(28,44),
			out1               => s_out1(28,44),
			out2               => s_out2(28,44),
			lock_lower_row_out => s_locks_lower_out(28,44),
			lock_lower_row_in  => s_locks_lower_in(28,44),
			in1                => s_in1(28,44),
			in2                => s_in2(28,44),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(44)
		);
	s_in1(28,44)            <= s_out1(29,44);
	s_in2(28,44)            <= s_out2(29,45);
	s_locks_lower_in(28,44) <= s_locks_lower_out(29,44);

		normal_cell_28_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,45),
			fetch              => s_fetch(28,45),
			data_in            => s_data_in(28,45),
			data_out           => s_data_out(28,45),
			out1               => s_out1(28,45),
			out2               => s_out2(28,45),
			lock_lower_row_out => s_locks_lower_out(28,45),
			lock_lower_row_in  => s_locks_lower_in(28,45),
			in1                => s_in1(28,45),
			in2                => s_in2(28,45),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(45)
		);
	s_in1(28,45)            <= s_out1(29,45);
	s_in2(28,45)            <= s_out2(29,46);
	s_locks_lower_in(28,45) <= s_locks_lower_out(29,45);

		normal_cell_28_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,46),
			fetch              => s_fetch(28,46),
			data_in            => s_data_in(28,46),
			data_out           => s_data_out(28,46),
			out1               => s_out1(28,46),
			out2               => s_out2(28,46),
			lock_lower_row_out => s_locks_lower_out(28,46),
			lock_lower_row_in  => s_locks_lower_in(28,46),
			in1                => s_in1(28,46),
			in2                => s_in2(28,46),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(46)
		);
	s_in1(28,46)            <= s_out1(29,46);
	s_in2(28,46)            <= s_out2(29,47);
	s_locks_lower_in(28,46) <= s_locks_lower_out(29,46);

		normal_cell_28_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,47),
			fetch              => s_fetch(28,47),
			data_in            => s_data_in(28,47),
			data_out           => s_data_out(28,47),
			out1               => s_out1(28,47),
			out2               => s_out2(28,47),
			lock_lower_row_out => s_locks_lower_out(28,47),
			lock_lower_row_in  => s_locks_lower_in(28,47),
			in1                => s_in1(28,47),
			in2                => s_in2(28,47),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(47)
		);
	s_in1(28,47)            <= s_out1(29,47);
	s_in2(28,47)            <= s_out2(29,48);
	s_locks_lower_in(28,47) <= s_locks_lower_out(29,47);

		normal_cell_28_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,48),
			fetch              => s_fetch(28,48),
			data_in            => s_data_in(28,48),
			data_out           => s_data_out(28,48),
			out1               => s_out1(28,48),
			out2               => s_out2(28,48),
			lock_lower_row_out => s_locks_lower_out(28,48),
			lock_lower_row_in  => s_locks_lower_in(28,48),
			in1                => s_in1(28,48),
			in2                => s_in2(28,48),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(48)
		);
	s_in1(28,48)            <= s_out1(29,48);
	s_in2(28,48)            <= s_out2(29,49);
	s_locks_lower_in(28,48) <= s_locks_lower_out(29,48);

		normal_cell_28_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,49),
			fetch              => s_fetch(28,49),
			data_in            => s_data_in(28,49),
			data_out           => s_data_out(28,49),
			out1               => s_out1(28,49),
			out2               => s_out2(28,49),
			lock_lower_row_out => s_locks_lower_out(28,49),
			lock_lower_row_in  => s_locks_lower_in(28,49),
			in1                => s_in1(28,49),
			in2                => s_in2(28,49),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(49)
		);
	s_in1(28,49)            <= s_out1(29,49);
	s_in2(28,49)            <= s_out2(29,50);
	s_locks_lower_in(28,49) <= s_locks_lower_out(29,49);

		normal_cell_28_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,50),
			fetch              => s_fetch(28,50),
			data_in            => s_data_in(28,50),
			data_out           => s_data_out(28,50),
			out1               => s_out1(28,50),
			out2               => s_out2(28,50),
			lock_lower_row_out => s_locks_lower_out(28,50),
			lock_lower_row_in  => s_locks_lower_in(28,50),
			in1                => s_in1(28,50),
			in2                => s_in2(28,50),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(50)
		);
	s_in1(28,50)            <= s_out1(29,50);
	s_in2(28,50)            <= s_out2(29,51);
	s_locks_lower_in(28,50) <= s_locks_lower_out(29,50);

		normal_cell_28_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,51),
			fetch              => s_fetch(28,51),
			data_in            => s_data_in(28,51),
			data_out           => s_data_out(28,51),
			out1               => s_out1(28,51),
			out2               => s_out2(28,51),
			lock_lower_row_out => s_locks_lower_out(28,51),
			lock_lower_row_in  => s_locks_lower_in(28,51),
			in1                => s_in1(28,51),
			in2                => s_in2(28,51),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(51)
		);
	s_in1(28,51)            <= s_out1(29,51);
	s_in2(28,51)            <= s_out2(29,52);
	s_locks_lower_in(28,51) <= s_locks_lower_out(29,51);

		normal_cell_28_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,52),
			fetch              => s_fetch(28,52),
			data_in            => s_data_in(28,52),
			data_out           => s_data_out(28,52),
			out1               => s_out1(28,52),
			out2               => s_out2(28,52),
			lock_lower_row_out => s_locks_lower_out(28,52),
			lock_lower_row_in  => s_locks_lower_in(28,52),
			in1                => s_in1(28,52),
			in2                => s_in2(28,52),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(52)
		);
	s_in1(28,52)            <= s_out1(29,52);
	s_in2(28,52)            <= s_out2(29,53);
	s_locks_lower_in(28,52) <= s_locks_lower_out(29,52);

		normal_cell_28_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,53),
			fetch              => s_fetch(28,53),
			data_in            => s_data_in(28,53),
			data_out           => s_data_out(28,53),
			out1               => s_out1(28,53),
			out2               => s_out2(28,53),
			lock_lower_row_out => s_locks_lower_out(28,53),
			lock_lower_row_in  => s_locks_lower_in(28,53),
			in1                => s_in1(28,53),
			in2                => s_in2(28,53),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(53)
		);
	s_in1(28,53)            <= s_out1(29,53);
	s_in2(28,53)            <= s_out2(29,54);
	s_locks_lower_in(28,53) <= s_locks_lower_out(29,53);

		normal_cell_28_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,54),
			fetch              => s_fetch(28,54),
			data_in            => s_data_in(28,54),
			data_out           => s_data_out(28,54),
			out1               => s_out1(28,54),
			out2               => s_out2(28,54),
			lock_lower_row_out => s_locks_lower_out(28,54),
			lock_lower_row_in  => s_locks_lower_in(28,54),
			in1                => s_in1(28,54),
			in2                => s_in2(28,54),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(54)
		);
	s_in1(28,54)            <= s_out1(29,54);
	s_in2(28,54)            <= s_out2(29,55);
	s_locks_lower_in(28,54) <= s_locks_lower_out(29,54);

		normal_cell_28_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,55),
			fetch              => s_fetch(28,55),
			data_in            => s_data_in(28,55),
			data_out           => s_data_out(28,55),
			out1               => s_out1(28,55),
			out2               => s_out2(28,55),
			lock_lower_row_out => s_locks_lower_out(28,55),
			lock_lower_row_in  => s_locks_lower_in(28,55),
			in1                => s_in1(28,55),
			in2                => s_in2(28,55),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(55)
		);
	s_in1(28,55)            <= s_out1(29,55);
	s_in2(28,55)            <= s_out2(29,56);
	s_locks_lower_in(28,55) <= s_locks_lower_out(29,55);

		normal_cell_28_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,56),
			fetch              => s_fetch(28,56),
			data_in            => s_data_in(28,56),
			data_out           => s_data_out(28,56),
			out1               => s_out1(28,56),
			out2               => s_out2(28,56),
			lock_lower_row_out => s_locks_lower_out(28,56),
			lock_lower_row_in  => s_locks_lower_in(28,56),
			in1                => s_in1(28,56),
			in2                => s_in2(28,56),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(56)
		);
	s_in1(28,56)            <= s_out1(29,56);
	s_in2(28,56)            <= s_out2(29,57);
	s_locks_lower_in(28,56) <= s_locks_lower_out(29,56);

		normal_cell_28_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,57),
			fetch              => s_fetch(28,57),
			data_in            => s_data_in(28,57),
			data_out           => s_data_out(28,57),
			out1               => s_out1(28,57),
			out2               => s_out2(28,57),
			lock_lower_row_out => s_locks_lower_out(28,57),
			lock_lower_row_in  => s_locks_lower_in(28,57),
			in1                => s_in1(28,57),
			in2                => s_in2(28,57),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(57)
		);
	s_in1(28,57)            <= s_out1(29,57);
	s_in2(28,57)            <= s_out2(29,58);
	s_locks_lower_in(28,57) <= s_locks_lower_out(29,57);

		normal_cell_28_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,58),
			fetch              => s_fetch(28,58),
			data_in            => s_data_in(28,58),
			data_out           => s_data_out(28,58),
			out1               => s_out1(28,58),
			out2               => s_out2(28,58),
			lock_lower_row_out => s_locks_lower_out(28,58),
			lock_lower_row_in  => s_locks_lower_in(28,58),
			in1                => s_in1(28,58),
			in2                => s_in2(28,58),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(58)
		);
	s_in1(28,58)            <= s_out1(29,58);
	s_in2(28,58)            <= s_out2(29,59);
	s_locks_lower_in(28,58) <= s_locks_lower_out(29,58);

		normal_cell_28_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,59),
			fetch              => s_fetch(28,59),
			data_in            => s_data_in(28,59),
			data_out           => s_data_out(28,59),
			out1               => s_out1(28,59),
			out2               => s_out2(28,59),
			lock_lower_row_out => s_locks_lower_out(28,59),
			lock_lower_row_in  => s_locks_lower_in(28,59),
			in1                => s_in1(28,59),
			in2                => s_in2(28,59),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(59)
		);
	s_in1(28,59)            <= s_out1(29,59);
	s_in2(28,59)            <= s_out2(29,60);
	s_locks_lower_in(28,59) <= s_locks_lower_out(29,59);

		last_col_cell_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(28,60),
			fetch              => s_fetch(28,60),
			data_in            => s_data_in(28,60),
			data_out           => s_data_out(28,60),
			out1               => s_out1(28,60),
			out2               => s_out2(28,60),
			lock_lower_row_out => s_locks_lower_out(28,60),
			lock_lower_row_in  => s_locks_lower_in(28,60),
			in1                => s_in1(28,60),
			in2                => (others => '0'),
			lock_row           => s_locks(28),
			piv_found          => s_piv_found,
			row_data           => s_row_data(28),
			col_data           => s_col_data(60)
		);
	s_in1(28,60)            <= s_out1(29,60);
	s_locks_lower_in(28,60) <= s_locks_lower_out(29,60);

		normal_cell_29_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,1),
			fetch              => s_fetch(29,1),
			data_in            => s_data_in(29,1),
			data_out           => s_data_out(29,1),
			out1               => s_out1(29,1),
			out2               => s_out2(29,1),
			lock_lower_row_out => s_locks_lower_out(29,1),
			lock_lower_row_in  => s_locks_lower_in(29,1),
			in1                => s_in1(29,1),
			in2                => s_in2(29,1),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(1)
		);
	s_in1(29,1)            <= s_out1(30,1);
	s_in2(29,1)            <= s_out2(30,2);
	s_locks_lower_in(29,1) <= s_locks_lower_out(30,1);

		normal_cell_29_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,2),
			fetch              => s_fetch(29,2),
			data_in            => s_data_in(29,2),
			data_out           => s_data_out(29,2),
			out1               => s_out1(29,2),
			out2               => s_out2(29,2),
			lock_lower_row_out => s_locks_lower_out(29,2),
			lock_lower_row_in  => s_locks_lower_in(29,2),
			in1                => s_in1(29,2),
			in2                => s_in2(29,2),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(2)
		);
	s_in1(29,2)            <= s_out1(30,2);
	s_in2(29,2)            <= s_out2(30,3);
	s_locks_lower_in(29,2) <= s_locks_lower_out(30,2);

		normal_cell_29_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,3),
			fetch              => s_fetch(29,3),
			data_in            => s_data_in(29,3),
			data_out           => s_data_out(29,3),
			out1               => s_out1(29,3),
			out2               => s_out2(29,3),
			lock_lower_row_out => s_locks_lower_out(29,3),
			lock_lower_row_in  => s_locks_lower_in(29,3),
			in1                => s_in1(29,3),
			in2                => s_in2(29,3),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(3)
		);
	s_in1(29,3)            <= s_out1(30,3);
	s_in2(29,3)            <= s_out2(30,4);
	s_locks_lower_in(29,3) <= s_locks_lower_out(30,3);

		normal_cell_29_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,4),
			fetch              => s_fetch(29,4),
			data_in            => s_data_in(29,4),
			data_out           => s_data_out(29,4),
			out1               => s_out1(29,4),
			out2               => s_out2(29,4),
			lock_lower_row_out => s_locks_lower_out(29,4),
			lock_lower_row_in  => s_locks_lower_in(29,4),
			in1                => s_in1(29,4),
			in2                => s_in2(29,4),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(4)
		);
	s_in1(29,4)            <= s_out1(30,4);
	s_in2(29,4)            <= s_out2(30,5);
	s_locks_lower_in(29,4) <= s_locks_lower_out(30,4);

		normal_cell_29_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,5),
			fetch              => s_fetch(29,5),
			data_in            => s_data_in(29,5),
			data_out           => s_data_out(29,5),
			out1               => s_out1(29,5),
			out2               => s_out2(29,5),
			lock_lower_row_out => s_locks_lower_out(29,5),
			lock_lower_row_in  => s_locks_lower_in(29,5),
			in1                => s_in1(29,5),
			in2                => s_in2(29,5),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(5)
		);
	s_in1(29,5)            <= s_out1(30,5);
	s_in2(29,5)            <= s_out2(30,6);
	s_locks_lower_in(29,5) <= s_locks_lower_out(30,5);

		normal_cell_29_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,6),
			fetch              => s_fetch(29,6),
			data_in            => s_data_in(29,6),
			data_out           => s_data_out(29,6),
			out1               => s_out1(29,6),
			out2               => s_out2(29,6),
			lock_lower_row_out => s_locks_lower_out(29,6),
			lock_lower_row_in  => s_locks_lower_in(29,6),
			in1                => s_in1(29,6),
			in2                => s_in2(29,6),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(6)
		);
	s_in1(29,6)            <= s_out1(30,6);
	s_in2(29,6)            <= s_out2(30,7);
	s_locks_lower_in(29,6) <= s_locks_lower_out(30,6);

		normal_cell_29_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,7),
			fetch              => s_fetch(29,7),
			data_in            => s_data_in(29,7),
			data_out           => s_data_out(29,7),
			out1               => s_out1(29,7),
			out2               => s_out2(29,7),
			lock_lower_row_out => s_locks_lower_out(29,7),
			lock_lower_row_in  => s_locks_lower_in(29,7),
			in1                => s_in1(29,7),
			in2                => s_in2(29,7),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(7)
		);
	s_in1(29,7)            <= s_out1(30,7);
	s_in2(29,7)            <= s_out2(30,8);
	s_locks_lower_in(29,7) <= s_locks_lower_out(30,7);

		normal_cell_29_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,8),
			fetch              => s_fetch(29,8),
			data_in            => s_data_in(29,8),
			data_out           => s_data_out(29,8),
			out1               => s_out1(29,8),
			out2               => s_out2(29,8),
			lock_lower_row_out => s_locks_lower_out(29,8),
			lock_lower_row_in  => s_locks_lower_in(29,8),
			in1                => s_in1(29,8),
			in2                => s_in2(29,8),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(8)
		);
	s_in1(29,8)            <= s_out1(30,8);
	s_in2(29,8)            <= s_out2(30,9);
	s_locks_lower_in(29,8) <= s_locks_lower_out(30,8);

		normal_cell_29_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,9),
			fetch              => s_fetch(29,9),
			data_in            => s_data_in(29,9),
			data_out           => s_data_out(29,9),
			out1               => s_out1(29,9),
			out2               => s_out2(29,9),
			lock_lower_row_out => s_locks_lower_out(29,9),
			lock_lower_row_in  => s_locks_lower_in(29,9),
			in1                => s_in1(29,9),
			in2                => s_in2(29,9),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(9)
		);
	s_in1(29,9)            <= s_out1(30,9);
	s_in2(29,9)            <= s_out2(30,10);
	s_locks_lower_in(29,9) <= s_locks_lower_out(30,9);

		normal_cell_29_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,10),
			fetch              => s_fetch(29,10),
			data_in            => s_data_in(29,10),
			data_out           => s_data_out(29,10),
			out1               => s_out1(29,10),
			out2               => s_out2(29,10),
			lock_lower_row_out => s_locks_lower_out(29,10),
			lock_lower_row_in  => s_locks_lower_in(29,10),
			in1                => s_in1(29,10),
			in2                => s_in2(29,10),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(10)
		);
	s_in1(29,10)            <= s_out1(30,10);
	s_in2(29,10)            <= s_out2(30,11);
	s_locks_lower_in(29,10) <= s_locks_lower_out(30,10);

		normal_cell_29_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,11),
			fetch              => s_fetch(29,11),
			data_in            => s_data_in(29,11),
			data_out           => s_data_out(29,11),
			out1               => s_out1(29,11),
			out2               => s_out2(29,11),
			lock_lower_row_out => s_locks_lower_out(29,11),
			lock_lower_row_in  => s_locks_lower_in(29,11),
			in1                => s_in1(29,11),
			in2                => s_in2(29,11),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(11)
		);
	s_in1(29,11)            <= s_out1(30,11);
	s_in2(29,11)            <= s_out2(30,12);
	s_locks_lower_in(29,11) <= s_locks_lower_out(30,11);

		normal_cell_29_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,12),
			fetch              => s_fetch(29,12),
			data_in            => s_data_in(29,12),
			data_out           => s_data_out(29,12),
			out1               => s_out1(29,12),
			out2               => s_out2(29,12),
			lock_lower_row_out => s_locks_lower_out(29,12),
			lock_lower_row_in  => s_locks_lower_in(29,12),
			in1                => s_in1(29,12),
			in2                => s_in2(29,12),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(12)
		);
	s_in1(29,12)            <= s_out1(30,12);
	s_in2(29,12)            <= s_out2(30,13);
	s_locks_lower_in(29,12) <= s_locks_lower_out(30,12);

		normal_cell_29_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,13),
			fetch              => s_fetch(29,13),
			data_in            => s_data_in(29,13),
			data_out           => s_data_out(29,13),
			out1               => s_out1(29,13),
			out2               => s_out2(29,13),
			lock_lower_row_out => s_locks_lower_out(29,13),
			lock_lower_row_in  => s_locks_lower_in(29,13),
			in1                => s_in1(29,13),
			in2                => s_in2(29,13),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(13)
		);
	s_in1(29,13)            <= s_out1(30,13);
	s_in2(29,13)            <= s_out2(30,14);
	s_locks_lower_in(29,13) <= s_locks_lower_out(30,13);

		normal_cell_29_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,14),
			fetch              => s_fetch(29,14),
			data_in            => s_data_in(29,14),
			data_out           => s_data_out(29,14),
			out1               => s_out1(29,14),
			out2               => s_out2(29,14),
			lock_lower_row_out => s_locks_lower_out(29,14),
			lock_lower_row_in  => s_locks_lower_in(29,14),
			in1                => s_in1(29,14),
			in2                => s_in2(29,14),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(14)
		);
	s_in1(29,14)            <= s_out1(30,14);
	s_in2(29,14)            <= s_out2(30,15);
	s_locks_lower_in(29,14) <= s_locks_lower_out(30,14);

		normal_cell_29_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,15),
			fetch              => s_fetch(29,15),
			data_in            => s_data_in(29,15),
			data_out           => s_data_out(29,15),
			out1               => s_out1(29,15),
			out2               => s_out2(29,15),
			lock_lower_row_out => s_locks_lower_out(29,15),
			lock_lower_row_in  => s_locks_lower_in(29,15),
			in1                => s_in1(29,15),
			in2                => s_in2(29,15),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(15)
		);
	s_in1(29,15)            <= s_out1(30,15);
	s_in2(29,15)            <= s_out2(30,16);
	s_locks_lower_in(29,15) <= s_locks_lower_out(30,15);

		normal_cell_29_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,16),
			fetch              => s_fetch(29,16),
			data_in            => s_data_in(29,16),
			data_out           => s_data_out(29,16),
			out1               => s_out1(29,16),
			out2               => s_out2(29,16),
			lock_lower_row_out => s_locks_lower_out(29,16),
			lock_lower_row_in  => s_locks_lower_in(29,16),
			in1                => s_in1(29,16),
			in2                => s_in2(29,16),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(16)
		);
	s_in1(29,16)            <= s_out1(30,16);
	s_in2(29,16)            <= s_out2(30,17);
	s_locks_lower_in(29,16) <= s_locks_lower_out(30,16);

		normal_cell_29_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,17),
			fetch              => s_fetch(29,17),
			data_in            => s_data_in(29,17),
			data_out           => s_data_out(29,17),
			out1               => s_out1(29,17),
			out2               => s_out2(29,17),
			lock_lower_row_out => s_locks_lower_out(29,17),
			lock_lower_row_in  => s_locks_lower_in(29,17),
			in1                => s_in1(29,17),
			in2                => s_in2(29,17),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(17)
		);
	s_in1(29,17)            <= s_out1(30,17);
	s_in2(29,17)            <= s_out2(30,18);
	s_locks_lower_in(29,17) <= s_locks_lower_out(30,17);

		normal_cell_29_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,18),
			fetch              => s_fetch(29,18),
			data_in            => s_data_in(29,18),
			data_out           => s_data_out(29,18),
			out1               => s_out1(29,18),
			out2               => s_out2(29,18),
			lock_lower_row_out => s_locks_lower_out(29,18),
			lock_lower_row_in  => s_locks_lower_in(29,18),
			in1                => s_in1(29,18),
			in2                => s_in2(29,18),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(18)
		);
	s_in1(29,18)            <= s_out1(30,18);
	s_in2(29,18)            <= s_out2(30,19);
	s_locks_lower_in(29,18) <= s_locks_lower_out(30,18);

		normal_cell_29_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,19),
			fetch              => s_fetch(29,19),
			data_in            => s_data_in(29,19),
			data_out           => s_data_out(29,19),
			out1               => s_out1(29,19),
			out2               => s_out2(29,19),
			lock_lower_row_out => s_locks_lower_out(29,19),
			lock_lower_row_in  => s_locks_lower_in(29,19),
			in1                => s_in1(29,19),
			in2                => s_in2(29,19),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(19)
		);
	s_in1(29,19)            <= s_out1(30,19);
	s_in2(29,19)            <= s_out2(30,20);
	s_locks_lower_in(29,19) <= s_locks_lower_out(30,19);

		normal_cell_29_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,20),
			fetch              => s_fetch(29,20),
			data_in            => s_data_in(29,20),
			data_out           => s_data_out(29,20),
			out1               => s_out1(29,20),
			out2               => s_out2(29,20),
			lock_lower_row_out => s_locks_lower_out(29,20),
			lock_lower_row_in  => s_locks_lower_in(29,20),
			in1                => s_in1(29,20),
			in2                => s_in2(29,20),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(20)
		);
	s_in1(29,20)            <= s_out1(30,20);
	s_in2(29,20)            <= s_out2(30,21);
	s_locks_lower_in(29,20) <= s_locks_lower_out(30,20);

		normal_cell_29_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,21),
			fetch              => s_fetch(29,21),
			data_in            => s_data_in(29,21),
			data_out           => s_data_out(29,21),
			out1               => s_out1(29,21),
			out2               => s_out2(29,21),
			lock_lower_row_out => s_locks_lower_out(29,21),
			lock_lower_row_in  => s_locks_lower_in(29,21),
			in1                => s_in1(29,21),
			in2                => s_in2(29,21),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(21)
		);
	s_in1(29,21)            <= s_out1(30,21);
	s_in2(29,21)            <= s_out2(30,22);
	s_locks_lower_in(29,21) <= s_locks_lower_out(30,21);

		normal_cell_29_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,22),
			fetch              => s_fetch(29,22),
			data_in            => s_data_in(29,22),
			data_out           => s_data_out(29,22),
			out1               => s_out1(29,22),
			out2               => s_out2(29,22),
			lock_lower_row_out => s_locks_lower_out(29,22),
			lock_lower_row_in  => s_locks_lower_in(29,22),
			in1                => s_in1(29,22),
			in2                => s_in2(29,22),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(22)
		);
	s_in1(29,22)            <= s_out1(30,22);
	s_in2(29,22)            <= s_out2(30,23);
	s_locks_lower_in(29,22) <= s_locks_lower_out(30,22);

		normal_cell_29_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,23),
			fetch              => s_fetch(29,23),
			data_in            => s_data_in(29,23),
			data_out           => s_data_out(29,23),
			out1               => s_out1(29,23),
			out2               => s_out2(29,23),
			lock_lower_row_out => s_locks_lower_out(29,23),
			lock_lower_row_in  => s_locks_lower_in(29,23),
			in1                => s_in1(29,23),
			in2                => s_in2(29,23),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(23)
		);
	s_in1(29,23)            <= s_out1(30,23);
	s_in2(29,23)            <= s_out2(30,24);
	s_locks_lower_in(29,23) <= s_locks_lower_out(30,23);

		normal_cell_29_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,24),
			fetch              => s_fetch(29,24),
			data_in            => s_data_in(29,24),
			data_out           => s_data_out(29,24),
			out1               => s_out1(29,24),
			out2               => s_out2(29,24),
			lock_lower_row_out => s_locks_lower_out(29,24),
			lock_lower_row_in  => s_locks_lower_in(29,24),
			in1                => s_in1(29,24),
			in2                => s_in2(29,24),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(24)
		);
	s_in1(29,24)            <= s_out1(30,24);
	s_in2(29,24)            <= s_out2(30,25);
	s_locks_lower_in(29,24) <= s_locks_lower_out(30,24);

		normal_cell_29_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,25),
			fetch              => s_fetch(29,25),
			data_in            => s_data_in(29,25),
			data_out           => s_data_out(29,25),
			out1               => s_out1(29,25),
			out2               => s_out2(29,25),
			lock_lower_row_out => s_locks_lower_out(29,25),
			lock_lower_row_in  => s_locks_lower_in(29,25),
			in1                => s_in1(29,25),
			in2                => s_in2(29,25),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(25)
		);
	s_in1(29,25)            <= s_out1(30,25);
	s_in2(29,25)            <= s_out2(30,26);
	s_locks_lower_in(29,25) <= s_locks_lower_out(30,25);

		normal_cell_29_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,26),
			fetch              => s_fetch(29,26),
			data_in            => s_data_in(29,26),
			data_out           => s_data_out(29,26),
			out1               => s_out1(29,26),
			out2               => s_out2(29,26),
			lock_lower_row_out => s_locks_lower_out(29,26),
			lock_lower_row_in  => s_locks_lower_in(29,26),
			in1                => s_in1(29,26),
			in2                => s_in2(29,26),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(26)
		);
	s_in1(29,26)            <= s_out1(30,26);
	s_in2(29,26)            <= s_out2(30,27);
	s_locks_lower_in(29,26) <= s_locks_lower_out(30,26);

		normal_cell_29_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,27),
			fetch              => s_fetch(29,27),
			data_in            => s_data_in(29,27),
			data_out           => s_data_out(29,27),
			out1               => s_out1(29,27),
			out2               => s_out2(29,27),
			lock_lower_row_out => s_locks_lower_out(29,27),
			lock_lower_row_in  => s_locks_lower_in(29,27),
			in1                => s_in1(29,27),
			in2                => s_in2(29,27),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(27)
		);
	s_in1(29,27)            <= s_out1(30,27);
	s_in2(29,27)            <= s_out2(30,28);
	s_locks_lower_in(29,27) <= s_locks_lower_out(30,27);

		normal_cell_29_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,28),
			fetch              => s_fetch(29,28),
			data_in            => s_data_in(29,28),
			data_out           => s_data_out(29,28),
			out1               => s_out1(29,28),
			out2               => s_out2(29,28),
			lock_lower_row_out => s_locks_lower_out(29,28),
			lock_lower_row_in  => s_locks_lower_in(29,28),
			in1                => s_in1(29,28),
			in2                => s_in2(29,28),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(28)
		);
	s_in1(29,28)            <= s_out1(30,28);
	s_in2(29,28)            <= s_out2(30,29);
	s_locks_lower_in(29,28) <= s_locks_lower_out(30,28);

		normal_cell_29_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,29),
			fetch              => s_fetch(29,29),
			data_in            => s_data_in(29,29),
			data_out           => s_data_out(29,29),
			out1               => s_out1(29,29),
			out2               => s_out2(29,29),
			lock_lower_row_out => s_locks_lower_out(29,29),
			lock_lower_row_in  => s_locks_lower_in(29,29),
			in1                => s_in1(29,29),
			in2                => s_in2(29,29),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(29)
		);
	s_in1(29,29)            <= s_out1(30,29);
	s_in2(29,29)            <= s_out2(30,30);
	s_locks_lower_in(29,29) <= s_locks_lower_out(30,29);

		normal_cell_29_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,30),
			fetch              => s_fetch(29,30),
			data_in            => s_data_in(29,30),
			data_out           => s_data_out(29,30),
			out1               => s_out1(29,30),
			out2               => s_out2(29,30),
			lock_lower_row_out => s_locks_lower_out(29,30),
			lock_lower_row_in  => s_locks_lower_in(29,30),
			in1                => s_in1(29,30),
			in2                => s_in2(29,30),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(30)
		);
	s_in1(29,30)            <= s_out1(30,30);
	s_in2(29,30)            <= s_out2(30,31);
	s_locks_lower_in(29,30) <= s_locks_lower_out(30,30);

		normal_cell_29_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,31),
			fetch              => s_fetch(29,31),
			data_in            => s_data_in(29,31),
			data_out           => s_data_out(29,31),
			out1               => s_out1(29,31),
			out2               => s_out2(29,31),
			lock_lower_row_out => s_locks_lower_out(29,31),
			lock_lower_row_in  => s_locks_lower_in(29,31),
			in1                => s_in1(29,31),
			in2                => s_in2(29,31),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(31)
		);
	s_in1(29,31)            <= s_out1(30,31);
	s_in2(29,31)            <= s_out2(30,32);
	s_locks_lower_in(29,31) <= s_locks_lower_out(30,31);

		normal_cell_29_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,32),
			fetch              => s_fetch(29,32),
			data_in            => s_data_in(29,32),
			data_out           => s_data_out(29,32),
			out1               => s_out1(29,32),
			out2               => s_out2(29,32),
			lock_lower_row_out => s_locks_lower_out(29,32),
			lock_lower_row_in  => s_locks_lower_in(29,32),
			in1                => s_in1(29,32),
			in2                => s_in2(29,32),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(32)
		);
	s_in1(29,32)            <= s_out1(30,32);
	s_in2(29,32)            <= s_out2(30,33);
	s_locks_lower_in(29,32) <= s_locks_lower_out(30,32);

		normal_cell_29_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,33),
			fetch              => s_fetch(29,33),
			data_in            => s_data_in(29,33),
			data_out           => s_data_out(29,33),
			out1               => s_out1(29,33),
			out2               => s_out2(29,33),
			lock_lower_row_out => s_locks_lower_out(29,33),
			lock_lower_row_in  => s_locks_lower_in(29,33),
			in1                => s_in1(29,33),
			in2                => s_in2(29,33),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(33)
		);
	s_in1(29,33)            <= s_out1(30,33);
	s_in2(29,33)            <= s_out2(30,34);
	s_locks_lower_in(29,33) <= s_locks_lower_out(30,33);

		normal_cell_29_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,34),
			fetch              => s_fetch(29,34),
			data_in            => s_data_in(29,34),
			data_out           => s_data_out(29,34),
			out1               => s_out1(29,34),
			out2               => s_out2(29,34),
			lock_lower_row_out => s_locks_lower_out(29,34),
			lock_lower_row_in  => s_locks_lower_in(29,34),
			in1                => s_in1(29,34),
			in2                => s_in2(29,34),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(34)
		);
	s_in1(29,34)            <= s_out1(30,34);
	s_in2(29,34)            <= s_out2(30,35);
	s_locks_lower_in(29,34) <= s_locks_lower_out(30,34);

		normal_cell_29_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,35),
			fetch              => s_fetch(29,35),
			data_in            => s_data_in(29,35),
			data_out           => s_data_out(29,35),
			out1               => s_out1(29,35),
			out2               => s_out2(29,35),
			lock_lower_row_out => s_locks_lower_out(29,35),
			lock_lower_row_in  => s_locks_lower_in(29,35),
			in1                => s_in1(29,35),
			in2                => s_in2(29,35),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(35)
		);
	s_in1(29,35)            <= s_out1(30,35);
	s_in2(29,35)            <= s_out2(30,36);
	s_locks_lower_in(29,35) <= s_locks_lower_out(30,35);

		normal_cell_29_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,36),
			fetch              => s_fetch(29,36),
			data_in            => s_data_in(29,36),
			data_out           => s_data_out(29,36),
			out1               => s_out1(29,36),
			out2               => s_out2(29,36),
			lock_lower_row_out => s_locks_lower_out(29,36),
			lock_lower_row_in  => s_locks_lower_in(29,36),
			in1                => s_in1(29,36),
			in2                => s_in2(29,36),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(36)
		);
	s_in1(29,36)            <= s_out1(30,36);
	s_in2(29,36)            <= s_out2(30,37);
	s_locks_lower_in(29,36) <= s_locks_lower_out(30,36);

		normal_cell_29_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,37),
			fetch              => s_fetch(29,37),
			data_in            => s_data_in(29,37),
			data_out           => s_data_out(29,37),
			out1               => s_out1(29,37),
			out2               => s_out2(29,37),
			lock_lower_row_out => s_locks_lower_out(29,37),
			lock_lower_row_in  => s_locks_lower_in(29,37),
			in1                => s_in1(29,37),
			in2                => s_in2(29,37),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(37)
		);
	s_in1(29,37)            <= s_out1(30,37);
	s_in2(29,37)            <= s_out2(30,38);
	s_locks_lower_in(29,37) <= s_locks_lower_out(30,37);

		normal_cell_29_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,38),
			fetch              => s_fetch(29,38),
			data_in            => s_data_in(29,38),
			data_out           => s_data_out(29,38),
			out1               => s_out1(29,38),
			out2               => s_out2(29,38),
			lock_lower_row_out => s_locks_lower_out(29,38),
			lock_lower_row_in  => s_locks_lower_in(29,38),
			in1                => s_in1(29,38),
			in2                => s_in2(29,38),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(38)
		);
	s_in1(29,38)            <= s_out1(30,38);
	s_in2(29,38)            <= s_out2(30,39);
	s_locks_lower_in(29,38) <= s_locks_lower_out(30,38);

		normal_cell_29_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,39),
			fetch              => s_fetch(29,39),
			data_in            => s_data_in(29,39),
			data_out           => s_data_out(29,39),
			out1               => s_out1(29,39),
			out2               => s_out2(29,39),
			lock_lower_row_out => s_locks_lower_out(29,39),
			lock_lower_row_in  => s_locks_lower_in(29,39),
			in1                => s_in1(29,39),
			in2                => s_in2(29,39),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(39)
		);
	s_in1(29,39)            <= s_out1(30,39);
	s_in2(29,39)            <= s_out2(30,40);
	s_locks_lower_in(29,39) <= s_locks_lower_out(30,39);

		normal_cell_29_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,40),
			fetch              => s_fetch(29,40),
			data_in            => s_data_in(29,40),
			data_out           => s_data_out(29,40),
			out1               => s_out1(29,40),
			out2               => s_out2(29,40),
			lock_lower_row_out => s_locks_lower_out(29,40),
			lock_lower_row_in  => s_locks_lower_in(29,40),
			in1                => s_in1(29,40),
			in2                => s_in2(29,40),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(40)
		);
	s_in1(29,40)            <= s_out1(30,40);
	s_in2(29,40)            <= s_out2(30,41);
	s_locks_lower_in(29,40) <= s_locks_lower_out(30,40);

		normal_cell_29_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,41),
			fetch              => s_fetch(29,41),
			data_in            => s_data_in(29,41),
			data_out           => s_data_out(29,41),
			out1               => s_out1(29,41),
			out2               => s_out2(29,41),
			lock_lower_row_out => s_locks_lower_out(29,41),
			lock_lower_row_in  => s_locks_lower_in(29,41),
			in1                => s_in1(29,41),
			in2                => s_in2(29,41),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(41)
		);
	s_in1(29,41)            <= s_out1(30,41);
	s_in2(29,41)            <= s_out2(30,42);
	s_locks_lower_in(29,41) <= s_locks_lower_out(30,41);

		normal_cell_29_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,42),
			fetch              => s_fetch(29,42),
			data_in            => s_data_in(29,42),
			data_out           => s_data_out(29,42),
			out1               => s_out1(29,42),
			out2               => s_out2(29,42),
			lock_lower_row_out => s_locks_lower_out(29,42),
			lock_lower_row_in  => s_locks_lower_in(29,42),
			in1                => s_in1(29,42),
			in2                => s_in2(29,42),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(42)
		);
	s_in1(29,42)            <= s_out1(30,42);
	s_in2(29,42)            <= s_out2(30,43);
	s_locks_lower_in(29,42) <= s_locks_lower_out(30,42);

		normal_cell_29_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,43),
			fetch              => s_fetch(29,43),
			data_in            => s_data_in(29,43),
			data_out           => s_data_out(29,43),
			out1               => s_out1(29,43),
			out2               => s_out2(29,43),
			lock_lower_row_out => s_locks_lower_out(29,43),
			lock_lower_row_in  => s_locks_lower_in(29,43),
			in1                => s_in1(29,43),
			in2                => s_in2(29,43),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(43)
		);
	s_in1(29,43)            <= s_out1(30,43);
	s_in2(29,43)            <= s_out2(30,44);
	s_locks_lower_in(29,43) <= s_locks_lower_out(30,43);

		normal_cell_29_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,44),
			fetch              => s_fetch(29,44),
			data_in            => s_data_in(29,44),
			data_out           => s_data_out(29,44),
			out1               => s_out1(29,44),
			out2               => s_out2(29,44),
			lock_lower_row_out => s_locks_lower_out(29,44),
			lock_lower_row_in  => s_locks_lower_in(29,44),
			in1                => s_in1(29,44),
			in2                => s_in2(29,44),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(44)
		);
	s_in1(29,44)            <= s_out1(30,44);
	s_in2(29,44)            <= s_out2(30,45);
	s_locks_lower_in(29,44) <= s_locks_lower_out(30,44);

		normal_cell_29_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,45),
			fetch              => s_fetch(29,45),
			data_in            => s_data_in(29,45),
			data_out           => s_data_out(29,45),
			out1               => s_out1(29,45),
			out2               => s_out2(29,45),
			lock_lower_row_out => s_locks_lower_out(29,45),
			lock_lower_row_in  => s_locks_lower_in(29,45),
			in1                => s_in1(29,45),
			in2                => s_in2(29,45),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(45)
		);
	s_in1(29,45)            <= s_out1(30,45);
	s_in2(29,45)            <= s_out2(30,46);
	s_locks_lower_in(29,45) <= s_locks_lower_out(30,45);

		normal_cell_29_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,46),
			fetch              => s_fetch(29,46),
			data_in            => s_data_in(29,46),
			data_out           => s_data_out(29,46),
			out1               => s_out1(29,46),
			out2               => s_out2(29,46),
			lock_lower_row_out => s_locks_lower_out(29,46),
			lock_lower_row_in  => s_locks_lower_in(29,46),
			in1                => s_in1(29,46),
			in2                => s_in2(29,46),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(46)
		);
	s_in1(29,46)            <= s_out1(30,46);
	s_in2(29,46)            <= s_out2(30,47);
	s_locks_lower_in(29,46) <= s_locks_lower_out(30,46);

		normal_cell_29_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,47),
			fetch              => s_fetch(29,47),
			data_in            => s_data_in(29,47),
			data_out           => s_data_out(29,47),
			out1               => s_out1(29,47),
			out2               => s_out2(29,47),
			lock_lower_row_out => s_locks_lower_out(29,47),
			lock_lower_row_in  => s_locks_lower_in(29,47),
			in1                => s_in1(29,47),
			in2                => s_in2(29,47),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(47)
		);
	s_in1(29,47)            <= s_out1(30,47);
	s_in2(29,47)            <= s_out2(30,48);
	s_locks_lower_in(29,47) <= s_locks_lower_out(30,47);

		normal_cell_29_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,48),
			fetch              => s_fetch(29,48),
			data_in            => s_data_in(29,48),
			data_out           => s_data_out(29,48),
			out1               => s_out1(29,48),
			out2               => s_out2(29,48),
			lock_lower_row_out => s_locks_lower_out(29,48),
			lock_lower_row_in  => s_locks_lower_in(29,48),
			in1                => s_in1(29,48),
			in2                => s_in2(29,48),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(48)
		);
	s_in1(29,48)            <= s_out1(30,48);
	s_in2(29,48)            <= s_out2(30,49);
	s_locks_lower_in(29,48) <= s_locks_lower_out(30,48);

		normal_cell_29_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,49),
			fetch              => s_fetch(29,49),
			data_in            => s_data_in(29,49),
			data_out           => s_data_out(29,49),
			out1               => s_out1(29,49),
			out2               => s_out2(29,49),
			lock_lower_row_out => s_locks_lower_out(29,49),
			lock_lower_row_in  => s_locks_lower_in(29,49),
			in1                => s_in1(29,49),
			in2                => s_in2(29,49),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(49)
		);
	s_in1(29,49)            <= s_out1(30,49);
	s_in2(29,49)            <= s_out2(30,50);
	s_locks_lower_in(29,49) <= s_locks_lower_out(30,49);

		normal_cell_29_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,50),
			fetch              => s_fetch(29,50),
			data_in            => s_data_in(29,50),
			data_out           => s_data_out(29,50),
			out1               => s_out1(29,50),
			out2               => s_out2(29,50),
			lock_lower_row_out => s_locks_lower_out(29,50),
			lock_lower_row_in  => s_locks_lower_in(29,50),
			in1                => s_in1(29,50),
			in2                => s_in2(29,50),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(50)
		);
	s_in1(29,50)            <= s_out1(30,50);
	s_in2(29,50)            <= s_out2(30,51);
	s_locks_lower_in(29,50) <= s_locks_lower_out(30,50);

		normal_cell_29_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,51),
			fetch              => s_fetch(29,51),
			data_in            => s_data_in(29,51),
			data_out           => s_data_out(29,51),
			out1               => s_out1(29,51),
			out2               => s_out2(29,51),
			lock_lower_row_out => s_locks_lower_out(29,51),
			lock_lower_row_in  => s_locks_lower_in(29,51),
			in1                => s_in1(29,51),
			in2                => s_in2(29,51),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(51)
		);
	s_in1(29,51)            <= s_out1(30,51);
	s_in2(29,51)            <= s_out2(30,52);
	s_locks_lower_in(29,51) <= s_locks_lower_out(30,51);

		normal_cell_29_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,52),
			fetch              => s_fetch(29,52),
			data_in            => s_data_in(29,52),
			data_out           => s_data_out(29,52),
			out1               => s_out1(29,52),
			out2               => s_out2(29,52),
			lock_lower_row_out => s_locks_lower_out(29,52),
			lock_lower_row_in  => s_locks_lower_in(29,52),
			in1                => s_in1(29,52),
			in2                => s_in2(29,52),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(52)
		);
	s_in1(29,52)            <= s_out1(30,52);
	s_in2(29,52)            <= s_out2(30,53);
	s_locks_lower_in(29,52) <= s_locks_lower_out(30,52);

		normal_cell_29_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,53),
			fetch              => s_fetch(29,53),
			data_in            => s_data_in(29,53),
			data_out           => s_data_out(29,53),
			out1               => s_out1(29,53),
			out2               => s_out2(29,53),
			lock_lower_row_out => s_locks_lower_out(29,53),
			lock_lower_row_in  => s_locks_lower_in(29,53),
			in1                => s_in1(29,53),
			in2                => s_in2(29,53),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(53)
		);
	s_in1(29,53)            <= s_out1(30,53);
	s_in2(29,53)            <= s_out2(30,54);
	s_locks_lower_in(29,53) <= s_locks_lower_out(30,53);

		normal_cell_29_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,54),
			fetch              => s_fetch(29,54),
			data_in            => s_data_in(29,54),
			data_out           => s_data_out(29,54),
			out1               => s_out1(29,54),
			out2               => s_out2(29,54),
			lock_lower_row_out => s_locks_lower_out(29,54),
			lock_lower_row_in  => s_locks_lower_in(29,54),
			in1                => s_in1(29,54),
			in2                => s_in2(29,54),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(54)
		);
	s_in1(29,54)            <= s_out1(30,54);
	s_in2(29,54)            <= s_out2(30,55);
	s_locks_lower_in(29,54) <= s_locks_lower_out(30,54);

		normal_cell_29_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,55),
			fetch              => s_fetch(29,55),
			data_in            => s_data_in(29,55),
			data_out           => s_data_out(29,55),
			out1               => s_out1(29,55),
			out2               => s_out2(29,55),
			lock_lower_row_out => s_locks_lower_out(29,55),
			lock_lower_row_in  => s_locks_lower_in(29,55),
			in1                => s_in1(29,55),
			in2                => s_in2(29,55),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(55)
		);
	s_in1(29,55)            <= s_out1(30,55);
	s_in2(29,55)            <= s_out2(30,56);
	s_locks_lower_in(29,55) <= s_locks_lower_out(30,55);

		normal_cell_29_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,56),
			fetch              => s_fetch(29,56),
			data_in            => s_data_in(29,56),
			data_out           => s_data_out(29,56),
			out1               => s_out1(29,56),
			out2               => s_out2(29,56),
			lock_lower_row_out => s_locks_lower_out(29,56),
			lock_lower_row_in  => s_locks_lower_in(29,56),
			in1                => s_in1(29,56),
			in2                => s_in2(29,56),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(56)
		);
	s_in1(29,56)            <= s_out1(30,56);
	s_in2(29,56)            <= s_out2(30,57);
	s_locks_lower_in(29,56) <= s_locks_lower_out(30,56);

		normal_cell_29_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,57),
			fetch              => s_fetch(29,57),
			data_in            => s_data_in(29,57),
			data_out           => s_data_out(29,57),
			out1               => s_out1(29,57),
			out2               => s_out2(29,57),
			lock_lower_row_out => s_locks_lower_out(29,57),
			lock_lower_row_in  => s_locks_lower_in(29,57),
			in1                => s_in1(29,57),
			in2                => s_in2(29,57),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(57)
		);
	s_in1(29,57)            <= s_out1(30,57);
	s_in2(29,57)            <= s_out2(30,58);
	s_locks_lower_in(29,57) <= s_locks_lower_out(30,57);

		normal_cell_29_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,58),
			fetch              => s_fetch(29,58),
			data_in            => s_data_in(29,58),
			data_out           => s_data_out(29,58),
			out1               => s_out1(29,58),
			out2               => s_out2(29,58),
			lock_lower_row_out => s_locks_lower_out(29,58),
			lock_lower_row_in  => s_locks_lower_in(29,58),
			in1                => s_in1(29,58),
			in2                => s_in2(29,58),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(58)
		);
	s_in1(29,58)            <= s_out1(30,58);
	s_in2(29,58)            <= s_out2(30,59);
	s_locks_lower_in(29,58) <= s_locks_lower_out(30,58);

		normal_cell_29_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,59),
			fetch              => s_fetch(29,59),
			data_in            => s_data_in(29,59),
			data_out           => s_data_out(29,59),
			out1               => s_out1(29,59),
			out2               => s_out2(29,59),
			lock_lower_row_out => s_locks_lower_out(29,59),
			lock_lower_row_in  => s_locks_lower_in(29,59),
			in1                => s_in1(29,59),
			in2                => s_in2(29,59),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(59)
		);
	s_in1(29,59)            <= s_out1(30,59);
	s_in2(29,59)            <= s_out2(30,60);
	s_locks_lower_in(29,59) <= s_locks_lower_out(30,59);

		last_col_cell_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(29,60),
			fetch              => s_fetch(29,60),
			data_in            => s_data_in(29,60),
			data_out           => s_data_out(29,60),
			out1               => s_out1(29,60),
			out2               => s_out2(29,60),
			lock_lower_row_out => s_locks_lower_out(29,60),
			lock_lower_row_in  => s_locks_lower_in(29,60),
			in1                => s_in1(29,60),
			in2                => (others => '0'),
			lock_row           => s_locks(29),
			piv_found          => s_piv_found,
			row_data           => s_row_data(29),
			col_data           => s_col_data(60)
		);
	s_in1(29,60)            <= s_out1(30,60);
	s_locks_lower_in(29,60) <= s_locks_lower_out(30,60);

		normal_cell_30_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,1),
			fetch              => s_fetch(30,1),
			data_in            => s_data_in(30,1),
			data_out           => s_data_out(30,1),
			out1               => s_out1(30,1),
			out2               => s_out2(30,1),
			lock_lower_row_out => s_locks_lower_out(30,1),
			lock_lower_row_in  => s_locks_lower_in(30,1),
			in1                => s_in1(30,1),
			in2                => s_in2(30,1),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(1)
		);
	s_in1(30,1)            <= s_out1(31,1);
	s_in2(30,1)            <= s_out2(31,2);
	s_locks_lower_in(30,1) <= s_locks_lower_out(31,1);

		normal_cell_30_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,2),
			fetch              => s_fetch(30,2),
			data_in            => s_data_in(30,2),
			data_out           => s_data_out(30,2),
			out1               => s_out1(30,2),
			out2               => s_out2(30,2),
			lock_lower_row_out => s_locks_lower_out(30,2),
			lock_lower_row_in  => s_locks_lower_in(30,2),
			in1                => s_in1(30,2),
			in2                => s_in2(30,2),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(2)
		);
	s_in1(30,2)            <= s_out1(31,2);
	s_in2(30,2)            <= s_out2(31,3);
	s_locks_lower_in(30,2) <= s_locks_lower_out(31,2);

		normal_cell_30_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,3),
			fetch              => s_fetch(30,3),
			data_in            => s_data_in(30,3),
			data_out           => s_data_out(30,3),
			out1               => s_out1(30,3),
			out2               => s_out2(30,3),
			lock_lower_row_out => s_locks_lower_out(30,3),
			lock_lower_row_in  => s_locks_lower_in(30,3),
			in1                => s_in1(30,3),
			in2                => s_in2(30,3),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(3)
		);
	s_in1(30,3)            <= s_out1(31,3);
	s_in2(30,3)            <= s_out2(31,4);
	s_locks_lower_in(30,3) <= s_locks_lower_out(31,3);

		normal_cell_30_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,4),
			fetch              => s_fetch(30,4),
			data_in            => s_data_in(30,4),
			data_out           => s_data_out(30,4),
			out1               => s_out1(30,4),
			out2               => s_out2(30,4),
			lock_lower_row_out => s_locks_lower_out(30,4),
			lock_lower_row_in  => s_locks_lower_in(30,4),
			in1                => s_in1(30,4),
			in2                => s_in2(30,4),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(4)
		);
	s_in1(30,4)            <= s_out1(31,4);
	s_in2(30,4)            <= s_out2(31,5);
	s_locks_lower_in(30,4) <= s_locks_lower_out(31,4);

		normal_cell_30_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,5),
			fetch              => s_fetch(30,5),
			data_in            => s_data_in(30,5),
			data_out           => s_data_out(30,5),
			out1               => s_out1(30,5),
			out2               => s_out2(30,5),
			lock_lower_row_out => s_locks_lower_out(30,5),
			lock_lower_row_in  => s_locks_lower_in(30,5),
			in1                => s_in1(30,5),
			in2                => s_in2(30,5),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(5)
		);
	s_in1(30,5)            <= s_out1(31,5);
	s_in2(30,5)            <= s_out2(31,6);
	s_locks_lower_in(30,5) <= s_locks_lower_out(31,5);

		normal_cell_30_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,6),
			fetch              => s_fetch(30,6),
			data_in            => s_data_in(30,6),
			data_out           => s_data_out(30,6),
			out1               => s_out1(30,6),
			out2               => s_out2(30,6),
			lock_lower_row_out => s_locks_lower_out(30,6),
			lock_lower_row_in  => s_locks_lower_in(30,6),
			in1                => s_in1(30,6),
			in2                => s_in2(30,6),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(6)
		);
	s_in1(30,6)            <= s_out1(31,6);
	s_in2(30,6)            <= s_out2(31,7);
	s_locks_lower_in(30,6) <= s_locks_lower_out(31,6);

		normal_cell_30_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,7),
			fetch              => s_fetch(30,7),
			data_in            => s_data_in(30,7),
			data_out           => s_data_out(30,7),
			out1               => s_out1(30,7),
			out2               => s_out2(30,7),
			lock_lower_row_out => s_locks_lower_out(30,7),
			lock_lower_row_in  => s_locks_lower_in(30,7),
			in1                => s_in1(30,7),
			in2                => s_in2(30,7),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(7)
		);
	s_in1(30,7)            <= s_out1(31,7);
	s_in2(30,7)            <= s_out2(31,8);
	s_locks_lower_in(30,7) <= s_locks_lower_out(31,7);

		normal_cell_30_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,8),
			fetch              => s_fetch(30,8),
			data_in            => s_data_in(30,8),
			data_out           => s_data_out(30,8),
			out1               => s_out1(30,8),
			out2               => s_out2(30,8),
			lock_lower_row_out => s_locks_lower_out(30,8),
			lock_lower_row_in  => s_locks_lower_in(30,8),
			in1                => s_in1(30,8),
			in2                => s_in2(30,8),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(8)
		);
	s_in1(30,8)            <= s_out1(31,8);
	s_in2(30,8)            <= s_out2(31,9);
	s_locks_lower_in(30,8) <= s_locks_lower_out(31,8);

		normal_cell_30_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,9),
			fetch              => s_fetch(30,9),
			data_in            => s_data_in(30,9),
			data_out           => s_data_out(30,9),
			out1               => s_out1(30,9),
			out2               => s_out2(30,9),
			lock_lower_row_out => s_locks_lower_out(30,9),
			lock_lower_row_in  => s_locks_lower_in(30,9),
			in1                => s_in1(30,9),
			in2                => s_in2(30,9),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(9)
		);
	s_in1(30,9)            <= s_out1(31,9);
	s_in2(30,9)            <= s_out2(31,10);
	s_locks_lower_in(30,9) <= s_locks_lower_out(31,9);

		normal_cell_30_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,10),
			fetch              => s_fetch(30,10),
			data_in            => s_data_in(30,10),
			data_out           => s_data_out(30,10),
			out1               => s_out1(30,10),
			out2               => s_out2(30,10),
			lock_lower_row_out => s_locks_lower_out(30,10),
			lock_lower_row_in  => s_locks_lower_in(30,10),
			in1                => s_in1(30,10),
			in2                => s_in2(30,10),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(10)
		);
	s_in1(30,10)            <= s_out1(31,10);
	s_in2(30,10)            <= s_out2(31,11);
	s_locks_lower_in(30,10) <= s_locks_lower_out(31,10);

		normal_cell_30_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,11),
			fetch              => s_fetch(30,11),
			data_in            => s_data_in(30,11),
			data_out           => s_data_out(30,11),
			out1               => s_out1(30,11),
			out2               => s_out2(30,11),
			lock_lower_row_out => s_locks_lower_out(30,11),
			lock_lower_row_in  => s_locks_lower_in(30,11),
			in1                => s_in1(30,11),
			in2                => s_in2(30,11),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(11)
		);
	s_in1(30,11)            <= s_out1(31,11);
	s_in2(30,11)            <= s_out2(31,12);
	s_locks_lower_in(30,11) <= s_locks_lower_out(31,11);

		normal_cell_30_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,12),
			fetch              => s_fetch(30,12),
			data_in            => s_data_in(30,12),
			data_out           => s_data_out(30,12),
			out1               => s_out1(30,12),
			out2               => s_out2(30,12),
			lock_lower_row_out => s_locks_lower_out(30,12),
			lock_lower_row_in  => s_locks_lower_in(30,12),
			in1                => s_in1(30,12),
			in2                => s_in2(30,12),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(12)
		);
	s_in1(30,12)            <= s_out1(31,12);
	s_in2(30,12)            <= s_out2(31,13);
	s_locks_lower_in(30,12) <= s_locks_lower_out(31,12);

		normal_cell_30_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,13),
			fetch              => s_fetch(30,13),
			data_in            => s_data_in(30,13),
			data_out           => s_data_out(30,13),
			out1               => s_out1(30,13),
			out2               => s_out2(30,13),
			lock_lower_row_out => s_locks_lower_out(30,13),
			lock_lower_row_in  => s_locks_lower_in(30,13),
			in1                => s_in1(30,13),
			in2                => s_in2(30,13),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(13)
		);
	s_in1(30,13)            <= s_out1(31,13);
	s_in2(30,13)            <= s_out2(31,14);
	s_locks_lower_in(30,13) <= s_locks_lower_out(31,13);

		normal_cell_30_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,14),
			fetch              => s_fetch(30,14),
			data_in            => s_data_in(30,14),
			data_out           => s_data_out(30,14),
			out1               => s_out1(30,14),
			out2               => s_out2(30,14),
			lock_lower_row_out => s_locks_lower_out(30,14),
			lock_lower_row_in  => s_locks_lower_in(30,14),
			in1                => s_in1(30,14),
			in2                => s_in2(30,14),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(14)
		);
	s_in1(30,14)            <= s_out1(31,14);
	s_in2(30,14)            <= s_out2(31,15);
	s_locks_lower_in(30,14) <= s_locks_lower_out(31,14);

		normal_cell_30_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,15),
			fetch              => s_fetch(30,15),
			data_in            => s_data_in(30,15),
			data_out           => s_data_out(30,15),
			out1               => s_out1(30,15),
			out2               => s_out2(30,15),
			lock_lower_row_out => s_locks_lower_out(30,15),
			lock_lower_row_in  => s_locks_lower_in(30,15),
			in1                => s_in1(30,15),
			in2                => s_in2(30,15),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(15)
		);
	s_in1(30,15)            <= s_out1(31,15);
	s_in2(30,15)            <= s_out2(31,16);
	s_locks_lower_in(30,15) <= s_locks_lower_out(31,15);

		normal_cell_30_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,16),
			fetch              => s_fetch(30,16),
			data_in            => s_data_in(30,16),
			data_out           => s_data_out(30,16),
			out1               => s_out1(30,16),
			out2               => s_out2(30,16),
			lock_lower_row_out => s_locks_lower_out(30,16),
			lock_lower_row_in  => s_locks_lower_in(30,16),
			in1                => s_in1(30,16),
			in2                => s_in2(30,16),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(16)
		);
	s_in1(30,16)            <= s_out1(31,16);
	s_in2(30,16)            <= s_out2(31,17);
	s_locks_lower_in(30,16) <= s_locks_lower_out(31,16);

		normal_cell_30_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,17),
			fetch              => s_fetch(30,17),
			data_in            => s_data_in(30,17),
			data_out           => s_data_out(30,17),
			out1               => s_out1(30,17),
			out2               => s_out2(30,17),
			lock_lower_row_out => s_locks_lower_out(30,17),
			lock_lower_row_in  => s_locks_lower_in(30,17),
			in1                => s_in1(30,17),
			in2                => s_in2(30,17),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(17)
		);
	s_in1(30,17)            <= s_out1(31,17);
	s_in2(30,17)            <= s_out2(31,18);
	s_locks_lower_in(30,17) <= s_locks_lower_out(31,17);

		normal_cell_30_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,18),
			fetch              => s_fetch(30,18),
			data_in            => s_data_in(30,18),
			data_out           => s_data_out(30,18),
			out1               => s_out1(30,18),
			out2               => s_out2(30,18),
			lock_lower_row_out => s_locks_lower_out(30,18),
			lock_lower_row_in  => s_locks_lower_in(30,18),
			in1                => s_in1(30,18),
			in2                => s_in2(30,18),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(18)
		);
	s_in1(30,18)            <= s_out1(31,18);
	s_in2(30,18)            <= s_out2(31,19);
	s_locks_lower_in(30,18) <= s_locks_lower_out(31,18);

		normal_cell_30_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,19),
			fetch              => s_fetch(30,19),
			data_in            => s_data_in(30,19),
			data_out           => s_data_out(30,19),
			out1               => s_out1(30,19),
			out2               => s_out2(30,19),
			lock_lower_row_out => s_locks_lower_out(30,19),
			lock_lower_row_in  => s_locks_lower_in(30,19),
			in1                => s_in1(30,19),
			in2                => s_in2(30,19),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(19)
		);
	s_in1(30,19)            <= s_out1(31,19);
	s_in2(30,19)            <= s_out2(31,20);
	s_locks_lower_in(30,19) <= s_locks_lower_out(31,19);

		normal_cell_30_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,20),
			fetch              => s_fetch(30,20),
			data_in            => s_data_in(30,20),
			data_out           => s_data_out(30,20),
			out1               => s_out1(30,20),
			out2               => s_out2(30,20),
			lock_lower_row_out => s_locks_lower_out(30,20),
			lock_lower_row_in  => s_locks_lower_in(30,20),
			in1                => s_in1(30,20),
			in2                => s_in2(30,20),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(20)
		);
	s_in1(30,20)            <= s_out1(31,20);
	s_in2(30,20)            <= s_out2(31,21);
	s_locks_lower_in(30,20) <= s_locks_lower_out(31,20);

		normal_cell_30_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,21),
			fetch              => s_fetch(30,21),
			data_in            => s_data_in(30,21),
			data_out           => s_data_out(30,21),
			out1               => s_out1(30,21),
			out2               => s_out2(30,21),
			lock_lower_row_out => s_locks_lower_out(30,21),
			lock_lower_row_in  => s_locks_lower_in(30,21),
			in1                => s_in1(30,21),
			in2                => s_in2(30,21),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(21)
		);
	s_in1(30,21)            <= s_out1(31,21);
	s_in2(30,21)            <= s_out2(31,22);
	s_locks_lower_in(30,21) <= s_locks_lower_out(31,21);

		normal_cell_30_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,22),
			fetch              => s_fetch(30,22),
			data_in            => s_data_in(30,22),
			data_out           => s_data_out(30,22),
			out1               => s_out1(30,22),
			out2               => s_out2(30,22),
			lock_lower_row_out => s_locks_lower_out(30,22),
			lock_lower_row_in  => s_locks_lower_in(30,22),
			in1                => s_in1(30,22),
			in2                => s_in2(30,22),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(22)
		);
	s_in1(30,22)            <= s_out1(31,22);
	s_in2(30,22)            <= s_out2(31,23);
	s_locks_lower_in(30,22) <= s_locks_lower_out(31,22);

		normal_cell_30_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,23),
			fetch              => s_fetch(30,23),
			data_in            => s_data_in(30,23),
			data_out           => s_data_out(30,23),
			out1               => s_out1(30,23),
			out2               => s_out2(30,23),
			lock_lower_row_out => s_locks_lower_out(30,23),
			lock_lower_row_in  => s_locks_lower_in(30,23),
			in1                => s_in1(30,23),
			in2                => s_in2(30,23),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(23)
		);
	s_in1(30,23)            <= s_out1(31,23);
	s_in2(30,23)            <= s_out2(31,24);
	s_locks_lower_in(30,23) <= s_locks_lower_out(31,23);

		normal_cell_30_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,24),
			fetch              => s_fetch(30,24),
			data_in            => s_data_in(30,24),
			data_out           => s_data_out(30,24),
			out1               => s_out1(30,24),
			out2               => s_out2(30,24),
			lock_lower_row_out => s_locks_lower_out(30,24),
			lock_lower_row_in  => s_locks_lower_in(30,24),
			in1                => s_in1(30,24),
			in2                => s_in2(30,24),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(24)
		);
	s_in1(30,24)            <= s_out1(31,24);
	s_in2(30,24)            <= s_out2(31,25);
	s_locks_lower_in(30,24) <= s_locks_lower_out(31,24);

		normal_cell_30_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,25),
			fetch              => s_fetch(30,25),
			data_in            => s_data_in(30,25),
			data_out           => s_data_out(30,25),
			out1               => s_out1(30,25),
			out2               => s_out2(30,25),
			lock_lower_row_out => s_locks_lower_out(30,25),
			lock_lower_row_in  => s_locks_lower_in(30,25),
			in1                => s_in1(30,25),
			in2                => s_in2(30,25),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(25)
		);
	s_in1(30,25)            <= s_out1(31,25);
	s_in2(30,25)            <= s_out2(31,26);
	s_locks_lower_in(30,25) <= s_locks_lower_out(31,25);

		normal_cell_30_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,26),
			fetch              => s_fetch(30,26),
			data_in            => s_data_in(30,26),
			data_out           => s_data_out(30,26),
			out1               => s_out1(30,26),
			out2               => s_out2(30,26),
			lock_lower_row_out => s_locks_lower_out(30,26),
			lock_lower_row_in  => s_locks_lower_in(30,26),
			in1                => s_in1(30,26),
			in2                => s_in2(30,26),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(26)
		);
	s_in1(30,26)            <= s_out1(31,26);
	s_in2(30,26)            <= s_out2(31,27);
	s_locks_lower_in(30,26) <= s_locks_lower_out(31,26);

		normal_cell_30_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,27),
			fetch              => s_fetch(30,27),
			data_in            => s_data_in(30,27),
			data_out           => s_data_out(30,27),
			out1               => s_out1(30,27),
			out2               => s_out2(30,27),
			lock_lower_row_out => s_locks_lower_out(30,27),
			lock_lower_row_in  => s_locks_lower_in(30,27),
			in1                => s_in1(30,27),
			in2                => s_in2(30,27),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(27)
		);
	s_in1(30,27)            <= s_out1(31,27);
	s_in2(30,27)            <= s_out2(31,28);
	s_locks_lower_in(30,27) <= s_locks_lower_out(31,27);

		normal_cell_30_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,28),
			fetch              => s_fetch(30,28),
			data_in            => s_data_in(30,28),
			data_out           => s_data_out(30,28),
			out1               => s_out1(30,28),
			out2               => s_out2(30,28),
			lock_lower_row_out => s_locks_lower_out(30,28),
			lock_lower_row_in  => s_locks_lower_in(30,28),
			in1                => s_in1(30,28),
			in2                => s_in2(30,28),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(28)
		);
	s_in1(30,28)            <= s_out1(31,28);
	s_in2(30,28)            <= s_out2(31,29);
	s_locks_lower_in(30,28) <= s_locks_lower_out(31,28);

		normal_cell_30_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,29),
			fetch              => s_fetch(30,29),
			data_in            => s_data_in(30,29),
			data_out           => s_data_out(30,29),
			out1               => s_out1(30,29),
			out2               => s_out2(30,29),
			lock_lower_row_out => s_locks_lower_out(30,29),
			lock_lower_row_in  => s_locks_lower_in(30,29),
			in1                => s_in1(30,29),
			in2                => s_in2(30,29),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(29)
		);
	s_in1(30,29)            <= s_out1(31,29);
	s_in2(30,29)            <= s_out2(31,30);
	s_locks_lower_in(30,29) <= s_locks_lower_out(31,29);

		normal_cell_30_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,30),
			fetch              => s_fetch(30,30),
			data_in            => s_data_in(30,30),
			data_out           => s_data_out(30,30),
			out1               => s_out1(30,30),
			out2               => s_out2(30,30),
			lock_lower_row_out => s_locks_lower_out(30,30),
			lock_lower_row_in  => s_locks_lower_in(30,30),
			in1                => s_in1(30,30),
			in2                => s_in2(30,30),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(30)
		);
	s_in1(30,30)            <= s_out1(31,30);
	s_in2(30,30)            <= s_out2(31,31);
	s_locks_lower_in(30,30) <= s_locks_lower_out(31,30);

		normal_cell_30_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,31),
			fetch              => s_fetch(30,31),
			data_in            => s_data_in(30,31),
			data_out           => s_data_out(30,31),
			out1               => s_out1(30,31),
			out2               => s_out2(30,31),
			lock_lower_row_out => s_locks_lower_out(30,31),
			lock_lower_row_in  => s_locks_lower_in(30,31),
			in1                => s_in1(30,31),
			in2                => s_in2(30,31),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(31)
		);
	s_in1(30,31)            <= s_out1(31,31);
	s_in2(30,31)            <= s_out2(31,32);
	s_locks_lower_in(30,31) <= s_locks_lower_out(31,31);

		normal_cell_30_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,32),
			fetch              => s_fetch(30,32),
			data_in            => s_data_in(30,32),
			data_out           => s_data_out(30,32),
			out1               => s_out1(30,32),
			out2               => s_out2(30,32),
			lock_lower_row_out => s_locks_lower_out(30,32),
			lock_lower_row_in  => s_locks_lower_in(30,32),
			in1                => s_in1(30,32),
			in2                => s_in2(30,32),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(32)
		);
	s_in1(30,32)            <= s_out1(31,32);
	s_in2(30,32)            <= s_out2(31,33);
	s_locks_lower_in(30,32) <= s_locks_lower_out(31,32);

		normal_cell_30_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,33),
			fetch              => s_fetch(30,33),
			data_in            => s_data_in(30,33),
			data_out           => s_data_out(30,33),
			out1               => s_out1(30,33),
			out2               => s_out2(30,33),
			lock_lower_row_out => s_locks_lower_out(30,33),
			lock_lower_row_in  => s_locks_lower_in(30,33),
			in1                => s_in1(30,33),
			in2                => s_in2(30,33),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(33)
		);
	s_in1(30,33)            <= s_out1(31,33);
	s_in2(30,33)            <= s_out2(31,34);
	s_locks_lower_in(30,33) <= s_locks_lower_out(31,33);

		normal_cell_30_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,34),
			fetch              => s_fetch(30,34),
			data_in            => s_data_in(30,34),
			data_out           => s_data_out(30,34),
			out1               => s_out1(30,34),
			out2               => s_out2(30,34),
			lock_lower_row_out => s_locks_lower_out(30,34),
			lock_lower_row_in  => s_locks_lower_in(30,34),
			in1                => s_in1(30,34),
			in2                => s_in2(30,34),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(34)
		);
	s_in1(30,34)            <= s_out1(31,34);
	s_in2(30,34)            <= s_out2(31,35);
	s_locks_lower_in(30,34) <= s_locks_lower_out(31,34);

		normal_cell_30_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,35),
			fetch              => s_fetch(30,35),
			data_in            => s_data_in(30,35),
			data_out           => s_data_out(30,35),
			out1               => s_out1(30,35),
			out2               => s_out2(30,35),
			lock_lower_row_out => s_locks_lower_out(30,35),
			lock_lower_row_in  => s_locks_lower_in(30,35),
			in1                => s_in1(30,35),
			in2                => s_in2(30,35),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(35)
		);
	s_in1(30,35)            <= s_out1(31,35);
	s_in2(30,35)            <= s_out2(31,36);
	s_locks_lower_in(30,35) <= s_locks_lower_out(31,35);

		normal_cell_30_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,36),
			fetch              => s_fetch(30,36),
			data_in            => s_data_in(30,36),
			data_out           => s_data_out(30,36),
			out1               => s_out1(30,36),
			out2               => s_out2(30,36),
			lock_lower_row_out => s_locks_lower_out(30,36),
			lock_lower_row_in  => s_locks_lower_in(30,36),
			in1                => s_in1(30,36),
			in2                => s_in2(30,36),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(36)
		);
	s_in1(30,36)            <= s_out1(31,36);
	s_in2(30,36)            <= s_out2(31,37);
	s_locks_lower_in(30,36) <= s_locks_lower_out(31,36);

		normal_cell_30_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,37),
			fetch              => s_fetch(30,37),
			data_in            => s_data_in(30,37),
			data_out           => s_data_out(30,37),
			out1               => s_out1(30,37),
			out2               => s_out2(30,37),
			lock_lower_row_out => s_locks_lower_out(30,37),
			lock_lower_row_in  => s_locks_lower_in(30,37),
			in1                => s_in1(30,37),
			in2                => s_in2(30,37),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(37)
		);
	s_in1(30,37)            <= s_out1(31,37);
	s_in2(30,37)            <= s_out2(31,38);
	s_locks_lower_in(30,37) <= s_locks_lower_out(31,37);

		normal_cell_30_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,38),
			fetch              => s_fetch(30,38),
			data_in            => s_data_in(30,38),
			data_out           => s_data_out(30,38),
			out1               => s_out1(30,38),
			out2               => s_out2(30,38),
			lock_lower_row_out => s_locks_lower_out(30,38),
			lock_lower_row_in  => s_locks_lower_in(30,38),
			in1                => s_in1(30,38),
			in2                => s_in2(30,38),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(38)
		);
	s_in1(30,38)            <= s_out1(31,38);
	s_in2(30,38)            <= s_out2(31,39);
	s_locks_lower_in(30,38) <= s_locks_lower_out(31,38);

		normal_cell_30_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,39),
			fetch              => s_fetch(30,39),
			data_in            => s_data_in(30,39),
			data_out           => s_data_out(30,39),
			out1               => s_out1(30,39),
			out2               => s_out2(30,39),
			lock_lower_row_out => s_locks_lower_out(30,39),
			lock_lower_row_in  => s_locks_lower_in(30,39),
			in1                => s_in1(30,39),
			in2                => s_in2(30,39),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(39)
		);
	s_in1(30,39)            <= s_out1(31,39);
	s_in2(30,39)            <= s_out2(31,40);
	s_locks_lower_in(30,39) <= s_locks_lower_out(31,39);

		normal_cell_30_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,40),
			fetch              => s_fetch(30,40),
			data_in            => s_data_in(30,40),
			data_out           => s_data_out(30,40),
			out1               => s_out1(30,40),
			out2               => s_out2(30,40),
			lock_lower_row_out => s_locks_lower_out(30,40),
			lock_lower_row_in  => s_locks_lower_in(30,40),
			in1                => s_in1(30,40),
			in2                => s_in2(30,40),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(40)
		);
	s_in1(30,40)            <= s_out1(31,40);
	s_in2(30,40)            <= s_out2(31,41);
	s_locks_lower_in(30,40) <= s_locks_lower_out(31,40);

		normal_cell_30_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,41),
			fetch              => s_fetch(30,41),
			data_in            => s_data_in(30,41),
			data_out           => s_data_out(30,41),
			out1               => s_out1(30,41),
			out2               => s_out2(30,41),
			lock_lower_row_out => s_locks_lower_out(30,41),
			lock_lower_row_in  => s_locks_lower_in(30,41),
			in1                => s_in1(30,41),
			in2                => s_in2(30,41),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(41)
		);
	s_in1(30,41)            <= s_out1(31,41);
	s_in2(30,41)            <= s_out2(31,42);
	s_locks_lower_in(30,41) <= s_locks_lower_out(31,41);

		normal_cell_30_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,42),
			fetch              => s_fetch(30,42),
			data_in            => s_data_in(30,42),
			data_out           => s_data_out(30,42),
			out1               => s_out1(30,42),
			out2               => s_out2(30,42),
			lock_lower_row_out => s_locks_lower_out(30,42),
			lock_lower_row_in  => s_locks_lower_in(30,42),
			in1                => s_in1(30,42),
			in2                => s_in2(30,42),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(42)
		);
	s_in1(30,42)            <= s_out1(31,42);
	s_in2(30,42)            <= s_out2(31,43);
	s_locks_lower_in(30,42) <= s_locks_lower_out(31,42);

		normal_cell_30_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,43),
			fetch              => s_fetch(30,43),
			data_in            => s_data_in(30,43),
			data_out           => s_data_out(30,43),
			out1               => s_out1(30,43),
			out2               => s_out2(30,43),
			lock_lower_row_out => s_locks_lower_out(30,43),
			lock_lower_row_in  => s_locks_lower_in(30,43),
			in1                => s_in1(30,43),
			in2                => s_in2(30,43),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(43)
		);
	s_in1(30,43)            <= s_out1(31,43);
	s_in2(30,43)            <= s_out2(31,44);
	s_locks_lower_in(30,43) <= s_locks_lower_out(31,43);

		normal_cell_30_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,44),
			fetch              => s_fetch(30,44),
			data_in            => s_data_in(30,44),
			data_out           => s_data_out(30,44),
			out1               => s_out1(30,44),
			out2               => s_out2(30,44),
			lock_lower_row_out => s_locks_lower_out(30,44),
			lock_lower_row_in  => s_locks_lower_in(30,44),
			in1                => s_in1(30,44),
			in2                => s_in2(30,44),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(44)
		);
	s_in1(30,44)            <= s_out1(31,44);
	s_in2(30,44)            <= s_out2(31,45);
	s_locks_lower_in(30,44) <= s_locks_lower_out(31,44);

		normal_cell_30_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,45),
			fetch              => s_fetch(30,45),
			data_in            => s_data_in(30,45),
			data_out           => s_data_out(30,45),
			out1               => s_out1(30,45),
			out2               => s_out2(30,45),
			lock_lower_row_out => s_locks_lower_out(30,45),
			lock_lower_row_in  => s_locks_lower_in(30,45),
			in1                => s_in1(30,45),
			in2                => s_in2(30,45),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(45)
		);
	s_in1(30,45)            <= s_out1(31,45);
	s_in2(30,45)            <= s_out2(31,46);
	s_locks_lower_in(30,45) <= s_locks_lower_out(31,45);

		normal_cell_30_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,46),
			fetch              => s_fetch(30,46),
			data_in            => s_data_in(30,46),
			data_out           => s_data_out(30,46),
			out1               => s_out1(30,46),
			out2               => s_out2(30,46),
			lock_lower_row_out => s_locks_lower_out(30,46),
			lock_lower_row_in  => s_locks_lower_in(30,46),
			in1                => s_in1(30,46),
			in2                => s_in2(30,46),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(46)
		);
	s_in1(30,46)            <= s_out1(31,46);
	s_in2(30,46)            <= s_out2(31,47);
	s_locks_lower_in(30,46) <= s_locks_lower_out(31,46);

		normal_cell_30_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,47),
			fetch              => s_fetch(30,47),
			data_in            => s_data_in(30,47),
			data_out           => s_data_out(30,47),
			out1               => s_out1(30,47),
			out2               => s_out2(30,47),
			lock_lower_row_out => s_locks_lower_out(30,47),
			lock_lower_row_in  => s_locks_lower_in(30,47),
			in1                => s_in1(30,47),
			in2                => s_in2(30,47),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(47)
		);
	s_in1(30,47)            <= s_out1(31,47);
	s_in2(30,47)            <= s_out2(31,48);
	s_locks_lower_in(30,47) <= s_locks_lower_out(31,47);

		normal_cell_30_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,48),
			fetch              => s_fetch(30,48),
			data_in            => s_data_in(30,48),
			data_out           => s_data_out(30,48),
			out1               => s_out1(30,48),
			out2               => s_out2(30,48),
			lock_lower_row_out => s_locks_lower_out(30,48),
			lock_lower_row_in  => s_locks_lower_in(30,48),
			in1                => s_in1(30,48),
			in2                => s_in2(30,48),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(48)
		);
	s_in1(30,48)            <= s_out1(31,48);
	s_in2(30,48)            <= s_out2(31,49);
	s_locks_lower_in(30,48) <= s_locks_lower_out(31,48);

		normal_cell_30_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,49),
			fetch              => s_fetch(30,49),
			data_in            => s_data_in(30,49),
			data_out           => s_data_out(30,49),
			out1               => s_out1(30,49),
			out2               => s_out2(30,49),
			lock_lower_row_out => s_locks_lower_out(30,49),
			lock_lower_row_in  => s_locks_lower_in(30,49),
			in1                => s_in1(30,49),
			in2                => s_in2(30,49),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(49)
		);
	s_in1(30,49)            <= s_out1(31,49);
	s_in2(30,49)            <= s_out2(31,50);
	s_locks_lower_in(30,49) <= s_locks_lower_out(31,49);

		normal_cell_30_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,50),
			fetch              => s_fetch(30,50),
			data_in            => s_data_in(30,50),
			data_out           => s_data_out(30,50),
			out1               => s_out1(30,50),
			out2               => s_out2(30,50),
			lock_lower_row_out => s_locks_lower_out(30,50),
			lock_lower_row_in  => s_locks_lower_in(30,50),
			in1                => s_in1(30,50),
			in2                => s_in2(30,50),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(50)
		);
	s_in1(30,50)            <= s_out1(31,50);
	s_in2(30,50)            <= s_out2(31,51);
	s_locks_lower_in(30,50) <= s_locks_lower_out(31,50);

		normal_cell_30_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,51),
			fetch              => s_fetch(30,51),
			data_in            => s_data_in(30,51),
			data_out           => s_data_out(30,51),
			out1               => s_out1(30,51),
			out2               => s_out2(30,51),
			lock_lower_row_out => s_locks_lower_out(30,51),
			lock_lower_row_in  => s_locks_lower_in(30,51),
			in1                => s_in1(30,51),
			in2                => s_in2(30,51),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(51)
		);
	s_in1(30,51)            <= s_out1(31,51);
	s_in2(30,51)            <= s_out2(31,52);
	s_locks_lower_in(30,51) <= s_locks_lower_out(31,51);

		normal_cell_30_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,52),
			fetch              => s_fetch(30,52),
			data_in            => s_data_in(30,52),
			data_out           => s_data_out(30,52),
			out1               => s_out1(30,52),
			out2               => s_out2(30,52),
			lock_lower_row_out => s_locks_lower_out(30,52),
			lock_lower_row_in  => s_locks_lower_in(30,52),
			in1                => s_in1(30,52),
			in2                => s_in2(30,52),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(52)
		);
	s_in1(30,52)            <= s_out1(31,52);
	s_in2(30,52)            <= s_out2(31,53);
	s_locks_lower_in(30,52) <= s_locks_lower_out(31,52);

		normal_cell_30_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,53),
			fetch              => s_fetch(30,53),
			data_in            => s_data_in(30,53),
			data_out           => s_data_out(30,53),
			out1               => s_out1(30,53),
			out2               => s_out2(30,53),
			lock_lower_row_out => s_locks_lower_out(30,53),
			lock_lower_row_in  => s_locks_lower_in(30,53),
			in1                => s_in1(30,53),
			in2                => s_in2(30,53),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(53)
		);
	s_in1(30,53)            <= s_out1(31,53);
	s_in2(30,53)            <= s_out2(31,54);
	s_locks_lower_in(30,53) <= s_locks_lower_out(31,53);

		normal_cell_30_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,54),
			fetch              => s_fetch(30,54),
			data_in            => s_data_in(30,54),
			data_out           => s_data_out(30,54),
			out1               => s_out1(30,54),
			out2               => s_out2(30,54),
			lock_lower_row_out => s_locks_lower_out(30,54),
			lock_lower_row_in  => s_locks_lower_in(30,54),
			in1                => s_in1(30,54),
			in2                => s_in2(30,54),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(54)
		);
	s_in1(30,54)            <= s_out1(31,54);
	s_in2(30,54)            <= s_out2(31,55);
	s_locks_lower_in(30,54) <= s_locks_lower_out(31,54);

		normal_cell_30_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,55),
			fetch              => s_fetch(30,55),
			data_in            => s_data_in(30,55),
			data_out           => s_data_out(30,55),
			out1               => s_out1(30,55),
			out2               => s_out2(30,55),
			lock_lower_row_out => s_locks_lower_out(30,55),
			lock_lower_row_in  => s_locks_lower_in(30,55),
			in1                => s_in1(30,55),
			in2                => s_in2(30,55),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(55)
		);
	s_in1(30,55)            <= s_out1(31,55);
	s_in2(30,55)            <= s_out2(31,56);
	s_locks_lower_in(30,55) <= s_locks_lower_out(31,55);

		normal_cell_30_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,56),
			fetch              => s_fetch(30,56),
			data_in            => s_data_in(30,56),
			data_out           => s_data_out(30,56),
			out1               => s_out1(30,56),
			out2               => s_out2(30,56),
			lock_lower_row_out => s_locks_lower_out(30,56),
			lock_lower_row_in  => s_locks_lower_in(30,56),
			in1                => s_in1(30,56),
			in2                => s_in2(30,56),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(56)
		);
	s_in1(30,56)            <= s_out1(31,56);
	s_in2(30,56)            <= s_out2(31,57);
	s_locks_lower_in(30,56) <= s_locks_lower_out(31,56);

		normal_cell_30_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,57),
			fetch              => s_fetch(30,57),
			data_in            => s_data_in(30,57),
			data_out           => s_data_out(30,57),
			out1               => s_out1(30,57),
			out2               => s_out2(30,57),
			lock_lower_row_out => s_locks_lower_out(30,57),
			lock_lower_row_in  => s_locks_lower_in(30,57),
			in1                => s_in1(30,57),
			in2                => s_in2(30,57),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(57)
		);
	s_in1(30,57)            <= s_out1(31,57);
	s_in2(30,57)            <= s_out2(31,58);
	s_locks_lower_in(30,57) <= s_locks_lower_out(31,57);

		normal_cell_30_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,58),
			fetch              => s_fetch(30,58),
			data_in            => s_data_in(30,58),
			data_out           => s_data_out(30,58),
			out1               => s_out1(30,58),
			out2               => s_out2(30,58),
			lock_lower_row_out => s_locks_lower_out(30,58),
			lock_lower_row_in  => s_locks_lower_in(30,58),
			in1                => s_in1(30,58),
			in2                => s_in2(30,58),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(58)
		);
	s_in1(30,58)            <= s_out1(31,58);
	s_in2(30,58)            <= s_out2(31,59);
	s_locks_lower_in(30,58) <= s_locks_lower_out(31,58);

		normal_cell_30_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,59),
			fetch              => s_fetch(30,59),
			data_in            => s_data_in(30,59),
			data_out           => s_data_out(30,59),
			out1               => s_out1(30,59),
			out2               => s_out2(30,59),
			lock_lower_row_out => s_locks_lower_out(30,59),
			lock_lower_row_in  => s_locks_lower_in(30,59),
			in1                => s_in1(30,59),
			in2                => s_in2(30,59),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(59)
		);
	s_in1(30,59)            <= s_out1(31,59);
	s_in2(30,59)            <= s_out2(31,60);
	s_locks_lower_in(30,59) <= s_locks_lower_out(31,59);

		last_col_cell_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(30,60),
			fetch              => s_fetch(30,60),
			data_in            => s_data_in(30,60),
			data_out           => s_data_out(30,60),
			out1               => s_out1(30,60),
			out2               => s_out2(30,60),
			lock_lower_row_out => s_locks_lower_out(30,60),
			lock_lower_row_in  => s_locks_lower_in(30,60),
			in1                => s_in1(30,60),
			in2                => (others => '0'),
			lock_row           => s_locks(30),
			piv_found          => s_piv_found,
			row_data           => s_row_data(30),
			col_data           => s_col_data(60)
		);
	s_in1(30,60)            <= s_out1(31,60);
	s_locks_lower_in(30,60) <= s_locks_lower_out(31,60);

		normal_cell_31_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,1),
			fetch              => s_fetch(31,1),
			data_in            => s_data_in(31,1),
			data_out           => s_data_out(31,1),
			out1               => s_out1(31,1),
			out2               => s_out2(31,1),
			lock_lower_row_out => s_locks_lower_out(31,1),
			lock_lower_row_in  => s_locks_lower_in(31,1),
			in1                => s_in1(31,1),
			in2                => s_in2(31,1),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(1)
		);
	s_in1(31,1)            <= s_out1(32,1);
	s_in2(31,1)            <= s_out2(32,2);
	s_locks_lower_in(31,1) <= s_locks_lower_out(32,1);

		normal_cell_31_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,2),
			fetch              => s_fetch(31,2),
			data_in            => s_data_in(31,2),
			data_out           => s_data_out(31,2),
			out1               => s_out1(31,2),
			out2               => s_out2(31,2),
			lock_lower_row_out => s_locks_lower_out(31,2),
			lock_lower_row_in  => s_locks_lower_in(31,2),
			in1                => s_in1(31,2),
			in2                => s_in2(31,2),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(2)
		);
	s_in1(31,2)            <= s_out1(32,2);
	s_in2(31,2)            <= s_out2(32,3);
	s_locks_lower_in(31,2) <= s_locks_lower_out(32,2);

		normal_cell_31_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,3),
			fetch              => s_fetch(31,3),
			data_in            => s_data_in(31,3),
			data_out           => s_data_out(31,3),
			out1               => s_out1(31,3),
			out2               => s_out2(31,3),
			lock_lower_row_out => s_locks_lower_out(31,3),
			lock_lower_row_in  => s_locks_lower_in(31,3),
			in1                => s_in1(31,3),
			in2                => s_in2(31,3),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(3)
		);
	s_in1(31,3)            <= s_out1(32,3);
	s_in2(31,3)            <= s_out2(32,4);
	s_locks_lower_in(31,3) <= s_locks_lower_out(32,3);

		normal_cell_31_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,4),
			fetch              => s_fetch(31,4),
			data_in            => s_data_in(31,4),
			data_out           => s_data_out(31,4),
			out1               => s_out1(31,4),
			out2               => s_out2(31,4),
			lock_lower_row_out => s_locks_lower_out(31,4),
			lock_lower_row_in  => s_locks_lower_in(31,4),
			in1                => s_in1(31,4),
			in2                => s_in2(31,4),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(4)
		);
	s_in1(31,4)            <= s_out1(32,4);
	s_in2(31,4)            <= s_out2(32,5);
	s_locks_lower_in(31,4) <= s_locks_lower_out(32,4);

		normal_cell_31_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,5),
			fetch              => s_fetch(31,5),
			data_in            => s_data_in(31,5),
			data_out           => s_data_out(31,5),
			out1               => s_out1(31,5),
			out2               => s_out2(31,5),
			lock_lower_row_out => s_locks_lower_out(31,5),
			lock_lower_row_in  => s_locks_lower_in(31,5),
			in1                => s_in1(31,5),
			in2                => s_in2(31,5),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(5)
		);
	s_in1(31,5)            <= s_out1(32,5);
	s_in2(31,5)            <= s_out2(32,6);
	s_locks_lower_in(31,5) <= s_locks_lower_out(32,5);

		normal_cell_31_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,6),
			fetch              => s_fetch(31,6),
			data_in            => s_data_in(31,6),
			data_out           => s_data_out(31,6),
			out1               => s_out1(31,6),
			out2               => s_out2(31,6),
			lock_lower_row_out => s_locks_lower_out(31,6),
			lock_lower_row_in  => s_locks_lower_in(31,6),
			in1                => s_in1(31,6),
			in2                => s_in2(31,6),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(6)
		);
	s_in1(31,6)            <= s_out1(32,6);
	s_in2(31,6)            <= s_out2(32,7);
	s_locks_lower_in(31,6) <= s_locks_lower_out(32,6);

		normal_cell_31_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,7),
			fetch              => s_fetch(31,7),
			data_in            => s_data_in(31,7),
			data_out           => s_data_out(31,7),
			out1               => s_out1(31,7),
			out2               => s_out2(31,7),
			lock_lower_row_out => s_locks_lower_out(31,7),
			lock_lower_row_in  => s_locks_lower_in(31,7),
			in1                => s_in1(31,7),
			in2                => s_in2(31,7),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(7)
		);
	s_in1(31,7)            <= s_out1(32,7);
	s_in2(31,7)            <= s_out2(32,8);
	s_locks_lower_in(31,7) <= s_locks_lower_out(32,7);

		normal_cell_31_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,8),
			fetch              => s_fetch(31,8),
			data_in            => s_data_in(31,8),
			data_out           => s_data_out(31,8),
			out1               => s_out1(31,8),
			out2               => s_out2(31,8),
			lock_lower_row_out => s_locks_lower_out(31,8),
			lock_lower_row_in  => s_locks_lower_in(31,8),
			in1                => s_in1(31,8),
			in2                => s_in2(31,8),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(8)
		);
	s_in1(31,8)            <= s_out1(32,8);
	s_in2(31,8)            <= s_out2(32,9);
	s_locks_lower_in(31,8) <= s_locks_lower_out(32,8);

		normal_cell_31_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,9),
			fetch              => s_fetch(31,9),
			data_in            => s_data_in(31,9),
			data_out           => s_data_out(31,9),
			out1               => s_out1(31,9),
			out2               => s_out2(31,9),
			lock_lower_row_out => s_locks_lower_out(31,9),
			lock_lower_row_in  => s_locks_lower_in(31,9),
			in1                => s_in1(31,9),
			in2                => s_in2(31,9),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(9)
		);
	s_in1(31,9)            <= s_out1(32,9);
	s_in2(31,9)            <= s_out2(32,10);
	s_locks_lower_in(31,9) <= s_locks_lower_out(32,9);

		normal_cell_31_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,10),
			fetch              => s_fetch(31,10),
			data_in            => s_data_in(31,10),
			data_out           => s_data_out(31,10),
			out1               => s_out1(31,10),
			out2               => s_out2(31,10),
			lock_lower_row_out => s_locks_lower_out(31,10),
			lock_lower_row_in  => s_locks_lower_in(31,10),
			in1                => s_in1(31,10),
			in2                => s_in2(31,10),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(10)
		);
	s_in1(31,10)            <= s_out1(32,10);
	s_in2(31,10)            <= s_out2(32,11);
	s_locks_lower_in(31,10) <= s_locks_lower_out(32,10);

		normal_cell_31_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,11),
			fetch              => s_fetch(31,11),
			data_in            => s_data_in(31,11),
			data_out           => s_data_out(31,11),
			out1               => s_out1(31,11),
			out2               => s_out2(31,11),
			lock_lower_row_out => s_locks_lower_out(31,11),
			lock_lower_row_in  => s_locks_lower_in(31,11),
			in1                => s_in1(31,11),
			in2                => s_in2(31,11),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(11)
		);
	s_in1(31,11)            <= s_out1(32,11);
	s_in2(31,11)            <= s_out2(32,12);
	s_locks_lower_in(31,11) <= s_locks_lower_out(32,11);

		normal_cell_31_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,12),
			fetch              => s_fetch(31,12),
			data_in            => s_data_in(31,12),
			data_out           => s_data_out(31,12),
			out1               => s_out1(31,12),
			out2               => s_out2(31,12),
			lock_lower_row_out => s_locks_lower_out(31,12),
			lock_lower_row_in  => s_locks_lower_in(31,12),
			in1                => s_in1(31,12),
			in2                => s_in2(31,12),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(12)
		);
	s_in1(31,12)            <= s_out1(32,12);
	s_in2(31,12)            <= s_out2(32,13);
	s_locks_lower_in(31,12) <= s_locks_lower_out(32,12);

		normal_cell_31_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,13),
			fetch              => s_fetch(31,13),
			data_in            => s_data_in(31,13),
			data_out           => s_data_out(31,13),
			out1               => s_out1(31,13),
			out2               => s_out2(31,13),
			lock_lower_row_out => s_locks_lower_out(31,13),
			lock_lower_row_in  => s_locks_lower_in(31,13),
			in1                => s_in1(31,13),
			in2                => s_in2(31,13),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(13)
		);
	s_in1(31,13)            <= s_out1(32,13);
	s_in2(31,13)            <= s_out2(32,14);
	s_locks_lower_in(31,13) <= s_locks_lower_out(32,13);

		normal_cell_31_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,14),
			fetch              => s_fetch(31,14),
			data_in            => s_data_in(31,14),
			data_out           => s_data_out(31,14),
			out1               => s_out1(31,14),
			out2               => s_out2(31,14),
			lock_lower_row_out => s_locks_lower_out(31,14),
			lock_lower_row_in  => s_locks_lower_in(31,14),
			in1                => s_in1(31,14),
			in2                => s_in2(31,14),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(14)
		);
	s_in1(31,14)            <= s_out1(32,14);
	s_in2(31,14)            <= s_out2(32,15);
	s_locks_lower_in(31,14) <= s_locks_lower_out(32,14);

		normal_cell_31_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,15),
			fetch              => s_fetch(31,15),
			data_in            => s_data_in(31,15),
			data_out           => s_data_out(31,15),
			out1               => s_out1(31,15),
			out2               => s_out2(31,15),
			lock_lower_row_out => s_locks_lower_out(31,15),
			lock_lower_row_in  => s_locks_lower_in(31,15),
			in1                => s_in1(31,15),
			in2                => s_in2(31,15),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(15)
		);
	s_in1(31,15)            <= s_out1(32,15);
	s_in2(31,15)            <= s_out2(32,16);
	s_locks_lower_in(31,15) <= s_locks_lower_out(32,15);

		normal_cell_31_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,16),
			fetch              => s_fetch(31,16),
			data_in            => s_data_in(31,16),
			data_out           => s_data_out(31,16),
			out1               => s_out1(31,16),
			out2               => s_out2(31,16),
			lock_lower_row_out => s_locks_lower_out(31,16),
			lock_lower_row_in  => s_locks_lower_in(31,16),
			in1                => s_in1(31,16),
			in2                => s_in2(31,16),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(16)
		);
	s_in1(31,16)            <= s_out1(32,16);
	s_in2(31,16)            <= s_out2(32,17);
	s_locks_lower_in(31,16) <= s_locks_lower_out(32,16);

		normal_cell_31_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,17),
			fetch              => s_fetch(31,17),
			data_in            => s_data_in(31,17),
			data_out           => s_data_out(31,17),
			out1               => s_out1(31,17),
			out2               => s_out2(31,17),
			lock_lower_row_out => s_locks_lower_out(31,17),
			lock_lower_row_in  => s_locks_lower_in(31,17),
			in1                => s_in1(31,17),
			in2                => s_in2(31,17),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(17)
		);
	s_in1(31,17)            <= s_out1(32,17);
	s_in2(31,17)            <= s_out2(32,18);
	s_locks_lower_in(31,17) <= s_locks_lower_out(32,17);

		normal_cell_31_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,18),
			fetch              => s_fetch(31,18),
			data_in            => s_data_in(31,18),
			data_out           => s_data_out(31,18),
			out1               => s_out1(31,18),
			out2               => s_out2(31,18),
			lock_lower_row_out => s_locks_lower_out(31,18),
			lock_lower_row_in  => s_locks_lower_in(31,18),
			in1                => s_in1(31,18),
			in2                => s_in2(31,18),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(18)
		);
	s_in1(31,18)            <= s_out1(32,18);
	s_in2(31,18)            <= s_out2(32,19);
	s_locks_lower_in(31,18) <= s_locks_lower_out(32,18);

		normal_cell_31_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,19),
			fetch              => s_fetch(31,19),
			data_in            => s_data_in(31,19),
			data_out           => s_data_out(31,19),
			out1               => s_out1(31,19),
			out2               => s_out2(31,19),
			lock_lower_row_out => s_locks_lower_out(31,19),
			lock_lower_row_in  => s_locks_lower_in(31,19),
			in1                => s_in1(31,19),
			in2                => s_in2(31,19),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(19)
		);
	s_in1(31,19)            <= s_out1(32,19);
	s_in2(31,19)            <= s_out2(32,20);
	s_locks_lower_in(31,19) <= s_locks_lower_out(32,19);

		normal_cell_31_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,20),
			fetch              => s_fetch(31,20),
			data_in            => s_data_in(31,20),
			data_out           => s_data_out(31,20),
			out1               => s_out1(31,20),
			out2               => s_out2(31,20),
			lock_lower_row_out => s_locks_lower_out(31,20),
			lock_lower_row_in  => s_locks_lower_in(31,20),
			in1                => s_in1(31,20),
			in2                => s_in2(31,20),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(20)
		);
	s_in1(31,20)            <= s_out1(32,20);
	s_in2(31,20)            <= s_out2(32,21);
	s_locks_lower_in(31,20) <= s_locks_lower_out(32,20);

		normal_cell_31_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,21),
			fetch              => s_fetch(31,21),
			data_in            => s_data_in(31,21),
			data_out           => s_data_out(31,21),
			out1               => s_out1(31,21),
			out2               => s_out2(31,21),
			lock_lower_row_out => s_locks_lower_out(31,21),
			lock_lower_row_in  => s_locks_lower_in(31,21),
			in1                => s_in1(31,21),
			in2                => s_in2(31,21),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(21)
		);
	s_in1(31,21)            <= s_out1(32,21);
	s_in2(31,21)            <= s_out2(32,22);
	s_locks_lower_in(31,21) <= s_locks_lower_out(32,21);

		normal_cell_31_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,22),
			fetch              => s_fetch(31,22),
			data_in            => s_data_in(31,22),
			data_out           => s_data_out(31,22),
			out1               => s_out1(31,22),
			out2               => s_out2(31,22),
			lock_lower_row_out => s_locks_lower_out(31,22),
			lock_lower_row_in  => s_locks_lower_in(31,22),
			in1                => s_in1(31,22),
			in2                => s_in2(31,22),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(22)
		);
	s_in1(31,22)            <= s_out1(32,22);
	s_in2(31,22)            <= s_out2(32,23);
	s_locks_lower_in(31,22) <= s_locks_lower_out(32,22);

		normal_cell_31_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,23),
			fetch              => s_fetch(31,23),
			data_in            => s_data_in(31,23),
			data_out           => s_data_out(31,23),
			out1               => s_out1(31,23),
			out2               => s_out2(31,23),
			lock_lower_row_out => s_locks_lower_out(31,23),
			lock_lower_row_in  => s_locks_lower_in(31,23),
			in1                => s_in1(31,23),
			in2                => s_in2(31,23),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(23)
		);
	s_in1(31,23)            <= s_out1(32,23);
	s_in2(31,23)            <= s_out2(32,24);
	s_locks_lower_in(31,23) <= s_locks_lower_out(32,23);

		normal_cell_31_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,24),
			fetch              => s_fetch(31,24),
			data_in            => s_data_in(31,24),
			data_out           => s_data_out(31,24),
			out1               => s_out1(31,24),
			out2               => s_out2(31,24),
			lock_lower_row_out => s_locks_lower_out(31,24),
			lock_lower_row_in  => s_locks_lower_in(31,24),
			in1                => s_in1(31,24),
			in2                => s_in2(31,24),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(24)
		);
	s_in1(31,24)            <= s_out1(32,24);
	s_in2(31,24)            <= s_out2(32,25);
	s_locks_lower_in(31,24) <= s_locks_lower_out(32,24);

		normal_cell_31_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,25),
			fetch              => s_fetch(31,25),
			data_in            => s_data_in(31,25),
			data_out           => s_data_out(31,25),
			out1               => s_out1(31,25),
			out2               => s_out2(31,25),
			lock_lower_row_out => s_locks_lower_out(31,25),
			lock_lower_row_in  => s_locks_lower_in(31,25),
			in1                => s_in1(31,25),
			in2                => s_in2(31,25),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(25)
		);
	s_in1(31,25)            <= s_out1(32,25);
	s_in2(31,25)            <= s_out2(32,26);
	s_locks_lower_in(31,25) <= s_locks_lower_out(32,25);

		normal_cell_31_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,26),
			fetch              => s_fetch(31,26),
			data_in            => s_data_in(31,26),
			data_out           => s_data_out(31,26),
			out1               => s_out1(31,26),
			out2               => s_out2(31,26),
			lock_lower_row_out => s_locks_lower_out(31,26),
			lock_lower_row_in  => s_locks_lower_in(31,26),
			in1                => s_in1(31,26),
			in2                => s_in2(31,26),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(26)
		);
	s_in1(31,26)            <= s_out1(32,26);
	s_in2(31,26)            <= s_out2(32,27);
	s_locks_lower_in(31,26) <= s_locks_lower_out(32,26);

		normal_cell_31_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,27),
			fetch              => s_fetch(31,27),
			data_in            => s_data_in(31,27),
			data_out           => s_data_out(31,27),
			out1               => s_out1(31,27),
			out2               => s_out2(31,27),
			lock_lower_row_out => s_locks_lower_out(31,27),
			lock_lower_row_in  => s_locks_lower_in(31,27),
			in1                => s_in1(31,27),
			in2                => s_in2(31,27),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(27)
		);
	s_in1(31,27)            <= s_out1(32,27);
	s_in2(31,27)            <= s_out2(32,28);
	s_locks_lower_in(31,27) <= s_locks_lower_out(32,27);

		normal_cell_31_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,28),
			fetch              => s_fetch(31,28),
			data_in            => s_data_in(31,28),
			data_out           => s_data_out(31,28),
			out1               => s_out1(31,28),
			out2               => s_out2(31,28),
			lock_lower_row_out => s_locks_lower_out(31,28),
			lock_lower_row_in  => s_locks_lower_in(31,28),
			in1                => s_in1(31,28),
			in2                => s_in2(31,28),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(28)
		);
	s_in1(31,28)            <= s_out1(32,28);
	s_in2(31,28)            <= s_out2(32,29);
	s_locks_lower_in(31,28) <= s_locks_lower_out(32,28);

		normal_cell_31_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,29),
			fetch              => s_fetch(31,29),
			data_in            => s_data_in(31,29),
			data_out           => s_data_out(31,29),
			out1               => s_out1(31,29),
			out2               => s_out2(31,29),
			lock_lower_row_out => s_locks_lower_out(31,29),
			lock_lower_row_in  => s_locks_lower_in(31,29),
			in1                => s_in1(31,29),
			in2                => s_in2(31,29),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(29)
		);
	s_in1(31,29)            <= s_out1(32,29);
	s_in2(31,29)            <= s_out2(32,30);
	s_locks_lower_in(31,29) <= s_locks_lower_out(32,29);

		normal_cell_31_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,30),
			fetch              => s_fetch(31,30),
			data_in            => s_data_in(31,30),
			data_out           => s_data_out(31,30),
			out1               => s_out1(31,30),
			out2               => s_out2(31,30),
			lock_lower_row_out => s_locks_lower_out(31,30),
			lock_lower_row_in  => s_locks_lower_in(31,30),
			in1                => s_in1(31,30),
			in2                => s_in2(31,30),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(30)
		);
	s_in1(31,30)            <= s_out1(32,30);
	s_in2(31,30)            <= s_out2(32,31);
	s_locks_lower_in(31,30) <= s_locks_lower_out(32,30);

		normal_cell_31_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,31),
			fetch              => s_fetch(31,31),
			data_in            => s_data_in(31,31),
			data_out           => s_data_out(31,31),
			out1               => s_out1(31,31),
			out2               => s_out2(31,31),
			lock_lower_row_out => s_locks_lower_out(31,31),
			lock_lower_row_in  => s_locks_lower_in(31,31),
			in1                => s_in1(31,31),
			in2                => s_in2(31,31),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(31)
		);
	s_in1(31,31)            <= s_out1(32,31);
	s_in2(31,31)            <= s_out2(32,32);
	s_locks_lower_in(31,31) <= s_locks_lower_out(32,31);

		normal_cell_31_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,32),
			fetch              => s_fetch(31,32),
			data_in            => s_data_in(31,32),
			data_out           => s_data_out(31,32),
			out1               => s_out1(31,32),
			out2               => s_out2(31,32),
			lock_lower_row_out => s_locks_lower_out(31,32),
			lock_lower_row_in  => s_locks_lower_in(31,32),
			in1                => s_in1(31,32),
			in2                => s_in2(31,32),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(32)
		);
	s_in1(31,32)            <= s_out1(32,32);
	s_in2(31,32)            <= s_out2(32,33);
	s_locks_lower_in(31,32) <= s_locks_lower_out(32,32);

		normal_cell_31_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,33),
			fetch              => s_fetch(31,33),
			data_in            => s_data_in(31,33),
			data_out           => s_data_out(31,33),
			out1               => s_out1(31,33),
			out2               => s_out2(31,33),
			lock_lower_row_out => s_locks_lower_out(31,33),
			lock_lower_row_in  => s_locks_lower_in(31,33),
			in1                => s_in1(31,33),
			in2                => s_in2(31,33),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(33)
		);
	s_in1(31,33)            <= s_out1(32,33);
	s_in2(31,33)            <= s_out2(32,34);
	s_locks_lower_in(31,33) <= s_locks_lower_out(32,33);

		normal_cell_31_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,34),
			fetch              => s_fetch(31,34),
			data_in            => s_data_in(31,34),
			data_out           => s_data_out(31,34),
			out1               => s_out1(31,34),
			out2               => s_out2(31,34),
			lock_lower_row_out => s_locks_lower_out(31,34),
			lock_lower_row_in  => s_locks_lower_in(31,34),
			in1                => s_in1(31,34),
			in2                => s_in2(31,34),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(34)
		);
	s_in1(31,34)            <= s_out1(32,34);
	s_in2(31,34)            <= s_out2(32,35);
	s_locks_lower_in(31,34) <= s_locks_lower_out(32,34);

		normal_cell_31_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,35),
			fetch              => s_fetch(31,35),
			data_in            => s_data_in(31,35),
			data_out           => s_data_out(31,35),
			out1               => s_out1(31,35),
			out2               => s_out2(31,35),
			lock_lower_row_out => s_locks_lower_out(31,35),
			lock_lower_row_in  => s_locks_lower_in(31,35),
			in1                => s_in1(31,35),
			in2                => s_in2(31,35),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(35)
		);
	s_in1(31,35)            <= s_out1(32,35);
	s_in2(31,35)            <= s_out2(32,36);
	s_locks_lower_in(31,35) <= s_locks_lower_out(32,35);

		normal_cell_31_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,36),
			fetch              => s_fetch(31,36),
			data_in            => s_data_in(31,36),
			data_out           => s_data_out(31,36),
			out1               => s_out1(31,36),
			out2               => s_out2(31,36),
			lock_lower_row_out => s_locks_lower_out(31,36),
			lock_lower_row_in  => s_locks_lower_in(31,36),
			in1                => s_in1(31,36),
			in2                => s_in2(31,36),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(36)
		);
	s_in1(31,36)            <= s_out1(32,36);
	s_in2(31,36)            <= s_out2(32,37);
	s_locks_lower_in(31,36) <= s_locks_lower_out(32,36);

		normal_cell_31_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,37),
			fetch              => s_fetch(31,37),
			data_in            => s_data_in(31,37),
			data_out           => s_data_out(31,37),
			out1               => s_out1(31,37),
			out2               => s_out2(31,37),
			lock_lower_row_out => s_locks_lower_out(31,37),
			lock_lower_row_in  => s_locks_lower_in(31,37),
			in1                => s_in1(31,37),
			in2                => s_in2(31,37),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(37)
		);
	s_in1(31,37)            <= s_out1(32,37);
	s_in2(31,37)            <= s_out2(32,38);
	s_locks_lower_in(31,37) <= s_locks_lower_out(32,37);

		normal_cell_31_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,38),
			fetch              => s_fetch(31,38),
			data_in            => s_data_in(31,38),
			data_out           => s_data_out(31,38),
			out1               => s_out1(31,38),
			out2               => s_out2(31,38),
			lock_lower_row_out => s_locks_lower_out(31,38),
			lock_lower_row_in  => s_locks_lower_in(31,38),
			in1                => s_in1(31,38),
			in2                => s_in2(31,38),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(38)
		);
	s_in1(31,38)            <= s_out1(32,38);
	s_in2(31,38)            <= s_out2(32,39);
	s_locks_lower_in(31,38) <= s_locks_lower_out(32,38);

		normal_cell_31_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,39),
			fetch              => s_fetch(31,39),
			data_in            => s_data_in(31,39),
			data_out           => s_data_out(31,39),
			out1               => s_out1(31,39),
			out2               => s_out2(31,39),
			lock_lower_row_out => s_locks_lower_out(31,39),
			lock_lower_row_in  => s_locks_lower_in(31,39),
			in1                => s_in1(31,39),
			in2                => s_in2(31,39),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(39)
		);
	s_in1(31,39)            <= s_out1(32,39);
	s_in2(31,39)            <= s_out2(32,40);
	s_locks_lower_in(31,39) <= s_locks_lower_out(32,39);

		normal_cell_31_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,40),
			fetch              => s_fetch(31,40),
			data_in            => s_data_in(31,40),
			data_out           => s_data_out(31,40),
			out1               => s_out1(31,40),
			out2               => s_out2(31,40),
			lock_lower_row_out => s_locks_lower_out(31,40),
			lock_lower_row_in  => s_locks_lower_in(31,40),
			in1                => s_in1(31,40),
			in2                => s_in2(31,40),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(40)
		);
	s_in1(31,40)            <= s_out1(32,40);
	s_in2(31,40)            <= s_out2(32,41);
	s_locks_lower_in(31,40) <= s_locks_lower_out(32,40);

		normal_cell_31_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,41),
			fetch              => s_fetch(31,41),
			data_in            => s_data_in(31,41),
			data_out           => s_data_out(31,41),
			out1               => s_out1(31,41),
			out2               => s_out2(31,41),
			lock_lower_row_out => s_locks_lower_out(31,41),
			lock_lower_row_in  => s_locks_lower_in(31,41),
			in1                => s_in1(31,41),
			in2                => s_in2(31,41),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(41)
		);
	s_in1(31,41)            <= s_out1(32,41);
	s_in2(31,41)            <= s_out2(32,42);
	s_locks_lower_in(31,41) <= s_locks_lower_out(32,41);

		normal_cell_31_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,42),
			fetch              => s_fetch(31,42),
			data_in            => s_data_in(31,42),
			data_out           => s_data_out(31,42),
			out1               => s_out1(31,42),
			out2               => s_out2(31,42),
			lock_lower_row_out => s_locks_lower_out(31,42),
			lock_lower_row_in  => s_locks_lower_in(31,42),
			in1                => s_in1(31,42),
			in2                => s_in2(31,42),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(42)
		);
	s_in1(31,42)            <= s_out1(32,42);
	s_in2(31,42)            <= s_out2(32,43);
	s_locks_lower_in(31,42) <= s_locks_lower_out(32,42);

		normal_cell_31_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,43),
			fetch              => s_fetch(31,43),
			data_in            => s_data_in(31,43),
			data_out           => s_data_out(31,43),
			out1               => s_out1(31,43),
			out2               => s_out2(31,43),
			lock_lower_row_out => s_locks_lower_out(31,43),
			lock_lower_row_in  => s_locks_lower_in(31,43),
			in1                => s_in1(31,43),
			in2                => s_in2(31,43),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(43)
		);
	s_in1(31,43)            <= s_out1(32,43);
	s_in2(31,43)            <= s_out2(32,44);
	s_locks_lower_in(31,43) <= s_locks_lower_out(32,43);

		normal_cell_31_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,44),
			fetch              => s_fetch(31,44),
			data_in            => s_data_in(31,44),
			data_out           => s_data_out(31,44),
			out1               => s_out1(31,44),
			out2               => s_out2(31,44),
			lock_lower_row_out => s_locks_lower_out(31,44),
			lock_lower_row_in  => s_locks_lower_in(31,44),
			in1                => s_in1(31,44),
			in2                => s_in2(31,44),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(44)
		);
	s_in1(31,44)            <= s_out1(32,44);
	s_in2(31,44)            <= s_out2(32,45);
	s_locks_lower_in(31,44) <= s_locks_lower_out(32,44);

		normal_cell_31_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,45),
			fetch              => s_fetch(31,45),
			data_in            => s_data_in(31,45),
			data_out           => s_data_out(31,45),
			out1               => s_out1(31,45),
			out2               => s_out2(31,45),
			lock_lower_row_out => s_locks_lower_out(31,45),
			lock_lower_row_in  => s_locks_lower_in(31,45),
			in1                => s_in1(31,45),
			in2                => s_in2(31,45),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(45)
		);
	s_in1(31,45)            <= s_out1(32,45);
	s_in2(31,45)            <= s_out2(32,46);
	s_locks_lower_in(31,45) <= s_locks_lower_out(32,45);

		normal_cell_31_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,46),
			fetch              => s_fetch(31,46),
			data_in            => s_data_in(31,46),
			data_out           => s_data_out(31,46),
			out1               => s_out1(31,46),
			out2               => s_out2(31,46),
			lock_lower_row_out => s_locks_lower_out(31,46),
			lock_lower_row_in  => s_locks_lower_in(31,46),
			in1                => s_in1(31,46),
			in2                => s_in2(31,46),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(46)
		);
	s_in1(31,46)            <= s_out1(32,46);
	s_in2(31,46)            <= s_out2(32,47);
	s_locks_lower_in(31,46) <= s_locks_lower_out(32,46);

		normal_cell_31_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,47),
			fetch              => s_fetch(31,47),
			data_in            => s_data_in(31,47),
			data_out           => s_data_out(31,47),
			out1               => s_out1(31,47),
			out2               => s_out2(31,47),
			lock_lower_row_out => s_locks_lower_out(31,47),
			lock_lower_row_in  => s_locks_lower_in(31,47),
			in1                => s_in1(31,47),
			in2                => s_in2(31,47),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(47)
		);
	s_in1(31,47)            <= s_out1(32,47);
	s_in2(31,47)            <= s_out2(32,48);
	s_locks_lower_in(31,47) <= s_locks_lower_out(32,47);

		normal_cell_31_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,48),
			fetch              => s_fetch(31,48),
			data_in            => s_data_in(31,48),
			data_out           => s_data_out(31,48),
			out1               => s_out1(31,48),
			out2               => s_out2(31,48),
			lock_lower_row_out => s_locks_lower_out(31,48),
			lock_lower_row_in  => s_locks_lower_in(31,48),
			in1                => s_in1(31,48),
			in2                => s_in2(31,48),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(48)
		);
	s_in1(31,48)            <= s_out1(32,48);
	s_in2(31,48)            <= s_out2(32,49);
	s_locks_lower_in(31,48) <= s_locks_lower_out(32,48);

		normal_cell_31_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,49),
			fetch              => s_fetch(31,49),
			data_in            => s_data_in(31,49),
			data_out           => s_data_out(31,49),
			out1               => s_out1(31,49),
			out2               => s_out2(31,49),
			lock_lower_row_out => s_locks_lower_out(31,49),
			lock_lower_row_in  => s_locks_lower_in(31,49),
			in1                => s_in1(31,49),
			in2                => s_in2(31,49),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(49)
		);
	s_in1(31,49)            <= s_out1(32,49);
	s_in2(31,49)            <= s_out2(32,50);
	s_locks_lower_in(31,49) <= s_locks_lower_out(32,49);

		normal_cell_31_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,50),
			fetch              => s_fetch(31,50),
			data_in            => s_data_in(31,50),
			data_out           => s_data_out(31,50),
			out1               => s_out1(31,50),
			out2               => s_out2(31,50),
			lock_lower_row_out => s_locks_lower_out(31,50),
			lock_lower_row_in  => s_locks_lower_in(31,50),
			in1                => s_in1(31,50),
			in2                => s_in2(31,50),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(50)
		);
	s_in1(31,50)            <= s_out1(32,50);
	s_in2(31,50)            <= s_out2(32,51);
	s_locks_lower_in(31,50) <= s_locks_lower_out(32,50);

		normal_cell_31_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,51),
			fetch              => s_fetch(31,51),
			data_in            => s_data_in(31,51),
			data_out           => s_data_out(31,51),
			out1               => s_out1(31,51),
			out2               => s_out2(31,51),
			lock_lower_row_out => s_locks_lower_out(31,51),
			lock_lower_row_in  => s_locks_lower_in(31,51),
			in1                => s_in1(31,51),
			in2                => s_in2(31,51),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(51)
		);
	s_in1(31,51)            <= s_out1(32,51);
	s_in2(31,51)            <= s_out2(32,52);
	s_locks_lower_in(31,51) <= s_locks_lower_out(32,51);

		normal_cell_31_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,52),
			fetch              => s_fetch(31,52),
			data_in            => s_data_in(31,52),
			data_out           => s_data_out(31,52),
			out1               => s_out1(31,52),
			out2               => s_out2(31,52),
			lock_lower_row_out => s_locks_lower_out(31,52),
			lock_lower_row_in  => s_locks_lower_in(31,52),
			in1                => s_in1(31,52),
			in2                => s_in2(31,52),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(52)
		);
	s_in1(31,52)            <= s_out1(32,52);
	s_in2(31,52)            <= s_out2(32,53);
	s_locks_lower_in(31,52) <= s_locks_lower_out(32,52);

		normal_cell_31_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,53),
			fetch              => s_fetch(31,53),
			data_in            => s_data_in(31,53),
			data_out           => s_data_out(31,53),
			out1               => s_out1(31,53),
			out2               => s_out2(31,53),
			lock_lower_row_out => s_locks_lower_out(31,53),
			lock_lower_row_in  => s_locks_lower_in(31,53),
			in1                => s_in1(31,53),
			in2                => s_in2(31,53),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(53)
		);
	s_in1(31,53)            <= s_out1(32,53);
	s_in2(31,53)            <= s_out2(32,54);
	s_locks_lower_in(31,53) <= s_locks_lower_out(32,53);

		normal_cell_31_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,54),
			fetch              => s_fetch(31,54),
			data_in            => s_data_in(31,54),
			data_out           => s_data_out(31,54),
			out1               => s_out1(31,54),
			out2               => s_out2(31,54),
			lock_lower_row_out => s_locks_lower_out(31,54),
			lock_lower_row_in  => s_locks_lower_in(31,54),
			in1                => s_in1(31,54),
			in2                => s_in2(31,54),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(54)
		);
	s_in1(31,54)            <= s_out1(32,54);
	s_in2(31,54)            <= s_out2(32,55);
	s_locks_lower_in(31,54) <= s_locks_lower_out(32,54);

		normal_cell_31_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,55),
			fetch              => s_fetch(31,55),
			data_in            => s_data_in(31,55),
			data_out           => s_data_out(31,55),
			out1               => s_out1(31,55),
			out2               => s_out2(31,55),
			lock_lower_row_out => s_locks_lower_out(31,55),
			lock_lower_row_in  => s_locks_lower_in(31,55),
			in1                => s_in1(31,55),
			in2                => s_in2(31,55),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(55)
		);
	s_in1(31,55)            <= s_out1(32,55);
	s_in2(31,55)            <= s_out2(32,56);
	s_locks_lower_in(31,55) <= s_locks_lower_out(32,55);

		normal_cell_31_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,56),
			fetch              => s_fetch(31,56),
			data_in            => s_data_in(31,56),
			data_out           => s_data_out(31,56),
			out1               => s_out1(31,56),
			out2               => s_out2(31,56),
			lock_lower_row_out => s_locks_lower_out(31,56),
			lock_lower_row_in  => s_locks_lower_in(31,56),
			in1                => s_in1(31,56),
			in2                => s_in2(31,56),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(56)
		);
	s_in1(31,56)            <= s_out1(32,56);
	s_in2(31,56)            <= s_out2(32,57);
	s_locks_lower_in(31,56) <= s_locks_lower_out(32,56);

		normal_cell_31_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,57),
			fetch              => s_fetch(31,57),
			data_in            => s_data_in(31,57),
			data_out           => s_data_out(31,57),
			out1               => s_out1(31,57),
			out2               => s_out2(31,57),
			lock_lower_row_out => s_locks_lower_out(31,57),
			lock_lower_row_in  => s_locks_lower_in(31,57),
			in1                => s_in1(31,57),
			in2                => s_in2(31,57),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(57)
		);
	s_in1(31,57)            <= s_out1(32,57);
	s_in2(31,57)            <= s_out2(32,58);
	s_locks_lower_in(31,57) <= s_locks_lower_out(32,57);

		normal_cell_31_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,58),
			fetch              => s_fetch(31,58),
			data_in            => s_data_in(31,58),
			data_out           => s_data_out(31,58),
			out1               => s_out1(31,58),
			out2               => s_out2(31,58),
			lock_lower_row_out => s_locks_lower_out(31,58),
			lock_lower_row_in  => s_locks_lower_in(31,58),
			in1                => s_in1(31,58),
			in2                => s_in2(31,58),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(58)
		);
	s_in1(31,58)            <= s_out1(32,58);
	s_in2(31,58)            <= s_out2(32,59);
	s_locks_lower_in(31,58) <= s_locks_lower_out(32,58);

		normal_cell_31_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,59),
			fetch              => s_fetch(31,59),
			data_in            => s_data_in(31,59),
			data_out           => s_data_out(31,59),
			out1               => s_out1(31,59),
			out2               => s_out2(31,59),
			lock_lower_row_out => s_locks_lower_out(31,59),
			lock_lower_row_in  => s_locks_lower_in(31,59),
			in1                => s_in1(31,59),
			in2                => s_in2(31,59),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(59)
		);
	s_in1(31,59)            <= s_out1(32,59);
	s_in2(31,59)            <= s_out2(32,60);
	s_locks_lower_in(31,59) <= s_locks_lower_out(32,59);

		last_col_cell_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(31,60),
			fetch              => s_fetch(31,60),
			data_in            => s_data_in(31,60),
			data_out           => s_data_out(31,60),
			out1               => s_out1(31,60),
			out2               => s_out2(31,60),
			lock_lower_row_out => s_locks_lower_out(31,60),
			lock_lower_row_in  => s_locks_lower_in(31,60),
			in1                => s_in1(31,60),
			in2                => (others => '0'),
			lock_row           => s_locks(31),
			piv_found          => s_piv_found,
			row_data           => s_row_data(31),
			col_data           => s_col_data(60)
		);
	s_in1(31,60)            <= s_out1(32,60);
	s_locks_lower_in(31,60) <= s_locks_lower_out(32,60);

		normal_cell_32_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,1),
			fetch              => s_fetch(32,1),
			data_in            => s_data_in(32,1),
			data_out           => s_data_out(32,1),
			out1               => s_out1(32,1),
			out2               => s_out2(32,1),
			lock_lower_row_out => s_locks_lower_out(32,1),
			lock_lower_row_in  => s_locks_lower_in(32,1),
			in1                => s_in1(32,1),
			in2                => s_in2(32,1),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(1)
		);
	s_in1(32,1)            <= s_out1(33,1);
	s_in2(32,1)            <= s_out2(33,2);
	s_locks_lower_in(32,1) <= s_locks_lower_out(33,1);

		normal_cell_32_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,2),
			fetch              => s_fetch(32,2),
			data_in            => s_data_in(32,2),
			data_out           => s_data_out(32,2),
			out1               => s_out1(32,2),
			out2               => s_out2(32,2),
			lock_lower_row_out => s_locks_lower_out(32,2),
			lock_lower_row_in  => s_locks_lower_in(32,2),
			in1                => s_in1(32,2),
			in2                => s_in2(32,2),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(2)
		);
	s_in1(32,2)            <= s_out1(33,2);
	s_in2(32,2)            <= s_out2(33,3);
	s_locks_lower_in(32,2) <= s_locks_lower_out(33,2);

		normal_cell_32_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,3),
			fetch              => s_fetch(32,3),
			data_in            => s_data_in(32,3),
			data_out           => s_data_out(32,3),
			out1               => s_out1(32,3),
			out2               => s_out2(32,3),
			lock_lower_row_out => s_locks_lower_out(32,3),
			lock_lower_row_in  => s_locks_lower_in(32,3),
			in1                => s_in1(32,3),
			in2                => s_in2(32,3),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(3)
		);
	s_in1(32,3)            <= s_out1(33,3);
	s_in2(32,3)            <= s_out2(33,4);
	s_locks_lower_in(32,3) <= s_locks_lower_out(33,3);

		normal_cell_32_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,4),
			fetch              => s_fetch(32,4),
			data_in            => s_data_in(32,4),
			data_out           => s_data_out(32,4),
			out1               => s_out1(32,4),
			out2               => s_out2(32,4),
			lock_lower_row_out => s_locks_lower_out(32,4),
			lock_lower_row_in  => s_locks_lower_in(32,4),
			in1                => s_in1(32,4),
			in2                => s_in2(32,4),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(4)
		);
	s_in1(32,4)            <= s_out1(33,4);
	s_in2(32,4)            <= s_out2(33,5);
	s_locks_lower_in(32,4) <= s_locks_lower_out(33,4);

		normal_cell_32_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,5),
			fetch              => s_fetch(32,5),
			data_in            => s_data_in(32,5),
			data_out           => s_data_out(32,5),
			out1               => s_out1(32,5),
			out2               => s_out2(32,5),
			lock_lower_row_out => s_locks_lower_out(32,5),
			lock_lower_row_in  => s_locks_lower_in(32,5),
			in1                => s_in1(32,5),
			in2                => s_in2(32,5),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(5)
		);
	s_in1(32,5)            <= s_out1(33,5);
	s_in2(32,5)            <= s_out2(33,6);
	s_locks_lower_in(32,5) <= s_locks_lower_out(33,5);

		normal_cell_32_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,6),
			fetch              => s_fetch(32,6),
			data_in            => s_data_in(32,6),
			data_out           => s_data_out(32,6),
			out1               => s_out1(32,6),
			out2               => s_out2(32,6),
			lock_lower_row_out => s_locks_lower_out(32,6),
			lock_lower_row_in  => s_locks_lower_in(32,6),
			in1                => s_in1(32,6),
			in2                => s_in2(32,6),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(6)
		);
	s_in1(32,6)            <= s_out1(33,6);
	s_in2(32,6)            <= s_out2(33,7);
	s_locks_lower_in(32,6) <= s_locks_lower_out(33,6);

		normal_cell_32_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,7),
			fetch              => s_fetch(32,7),
			data_in            => s_data_in(32,7),
			data_out           => s_data_out(32,7),
			out1               => s_out1(32,7),
			out2               => s_out2(32,7),
			lock_lower_row_out => s_locks_lower_out(32,7),
			lock_lower_row_in  => s_locks_lower_in(32,7),
			in1                => s_in1(32,7),
			in2                => s_in2(32,7),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(7)
		);
	s_in1(32,7)            <= s_out1(33,7);
	s_in2(32,7)            <= s_out2(33,8);
	s_locks_lower_in(32,7) <= s_locks_lower_out(33,7);

		normal_cell_32_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,8),
			fetch              => s_fetch(32,8),
			data_in            => s_data_in(32,8),
			data_out           => s_data_out(32,8),
			out1               => s_out1(32,8),
			out2               => s_out2(32,8),
			lock_lower_row_out => s_locks_lower_out(32,8),
			lock_lower_row_in  => s_locks_lower_in(32,8),
			in1                => s_in1(32,8),
			in2                => s_in2(32,8),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(8)
		);
	s_in1(32,8)            <= s_out1(33,8);
	s_in2(32,8)            <= s_out2(33,9);
	s_locks_lower_in(32,8) <= s_locks_lower_out(33,8);

		normal_cell_32_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,9),
			fetch              => s_fetch(32,9),
			data_in            => s_data_in(32,9),
			data_out           => s_data_out(32,9),
			out1               => s_out1(32,9),
			out2               => s_out2(32,9),
			lock_lower_row_out => s_locks_lower_out(32,9),
			lock_lower_row_in  => s_locks_lower_in(32,9),
			in1                => s_in1(32,9),
			in2                => s_in2(32,9),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(9)
		);
	s_in1(32,9)            <= s_out1(33,9);
	s_in2(32,9)            <= s_out2(33,10);
	s_locks_lower_in(32,9) <= s_locks_lower_out(33,9);

		normal_cell_32_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,10),
			fetch              => s_fetch(32,10),
			data_in            => s_data_in(32,10),
			data_out           => s_data_out(32,10),
			out1               => s_out1(32,10),
			out2               => s_out2(32,10),
			lock_lower_row_out => s_locks_lower_out(32,10),
			lock_lower_row_in  => s_locks_lower_in(32,10),
			in1                => s_in1(32,10),
			in2                => s_in2(32,10),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(10)
		);
	s_in1(32,10)            <= s_out1(33,10);
	s_in2(32,10)            <= s_out2(33,11);
	s_locks_lower_in(32,10) <= s_locks_lower_out(33,10);

		normal_cell_32_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,11),
			fetch              => s_fetch(32,11),
			data_in            => s_data_in(32,11),
			data_out           => s_data_out(32,11),
			out1               => s_out1(32,11),
			out2               => s_out2(32,11),
			lock_lower_row_out => s_locks_lower_out(32,11),
			lock_lower_row_in  => s_locks_lower_in(32,11),
			in1                => s_in1(32,11),
			in2                => s_in2(32,11),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(11)
		);
	s_in1(32,11)            <= s_out1(33,11);
	s_in2(32,11)            <= s_out2(33,12);
	s_locks_lower_in(32,11) <= s_locks_lower_out(33,11);

		normal_cell_32_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,12),
			fetch              => s_fetch(32,12),
			data_in            => s_data_in(32,12),
			data_out           => s_data_out(32,12),
			out1               => s_out1(32,12),
			out2               => s_out2(32,12),
			lock_lower_row_out => s_locks_lower_out(32,12),
			lock_lower_row_in  => s_locks_lower_in(32,12),
			in1                => s_in1(32,12),
			in2                => s_in2(32,12),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(12)
		);
	s_in1(32,12)            <= s_out1(33,12);
	s_in2(32,12)            <= s_out2(33,13);
	s_locks_lower_in(32,12) <= s_locks_lower_out(33,12);

		normal_cell_32_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,13),
			fetch              => s_fetch(32,13),
			data_in            => s_data_in(32,13),
			data_out           => s_data_out(32,13),
			out1               => s_out1(32,13),
			out2               => s_out2(32,13),
			lock_lower_row_out => s_locks_lower_out(32,13),
			lock_lower_row_in  => s_locks_lower_in(32,13),
			in1                => s_in1(32,13),
			in2                => s_in2(32,13),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(13)
		);
	s_in1(32,13)            <= s_out1(33,13);
	s_in2(32,13)            <= s_out2(33,14);
	s_locks_lower_in(32,13) <= s_locks_lower_out(33,13);

		normal_cell_32_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,14),
			fetch              => s_fetch(32,14),
			data_in            => s_data_in(32,14),
			data_out           => s_data_out(32,14),
			out1               => s_out1(32,14),
			out2               => s_out2(32,14),
			lock_lower_row_out => s_locks_lower_out(32,14),
			lock_lower_row_in  => s_locks_lower_in(32,14),
			in1                => s_in1(32,14),
			in2                => s_in2(32,14),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(14)
		);
	s_in1(32,14)            <= s_out1(33,14);
	s_in2(32,14)            <= s_out2(33,15);
	s_locks_lower_in(32,14) <= s_locks_lower_out(33,14);

		normal_cell_32_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,15),
			fetch              => s_fetch(32,15),
			data_in            => s_data_in(32,15),
			data_out           => s_data_out(32,15),
			out1               => s_out1(32,15),
			out2               => s_out2(32,15),
			lock_lower_row_out => s_locks_lower_out(32,15),
			lock_lower_row_in  => s_locks_lower_in(32,15),
			in1                => s_in1(32,15),
			in2                => s_in2(32,15),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(15)
		);
	s_in1(32,15)            <= s_out1(33,15);
	s_in2(32,15)            <= s_out2(33,16);
	s_locks_lower_in(32,15) <= s_locks_lower_out(33,15);

		normal_cell_32_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,16),
			fetch              => s_fetch(32,16),
			data_in            => s_data_in(32,16),
			data_out           => s_data_out(32,16),
			out1               => s_out1(32,16),
			out2               => s_out2(32,16),
			lock_lower_row_out => s_locks_lower_out(32,16),
			lock_lower_row_in  => s_locks_lower_in(32,16),
			in1                => s_in1(32,16),
			in2                => s_in2(32,16),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(16)
		);
	s_in1(32,16)            <= s_out1(33,16);
	s_in2(32,16)            <= s_out2(33,17);
	s_locks_lower_in(32,16) <= s_locks_lower_out(33,16);

		normal_cell_32_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,17),
			fetch              => s_fetch(32,17),
			data_in            => s_data_in(32,17),
			data_out           => s_data_out(32,17),
			out1               => s_out1(32,17),
			out2               => s_out2(32,17),
			lock_lower_row_out => s_locks_lower_out(32,17),
			lock_lower_row_in  => s_locks_lower_in(32,17),
			in1                => s_in1(32,17),
			in2                => s_in2(32,17),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(17)
		);
	s_in1(32,17)            <= s_out1(33,17);
	s_in2(32,17)            <= s_out2(33,18);
	s_locks_lower_in(32,17) <= s_locks_lower_out(33,17);

		normal_cell_32_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,18),
			fetch              => s_fetch(32,18),
			data_in            => s_data_in(32,18),
			data_out           => s_data_out(32,18),
			out1               => s_out1(32,18),
			out2               => s_out2(32,18),
			lock_lower_row_out => s_locks_lower_out(32,18),
			lock_lower_row_in  => s_locks_lower_in(32,18),
			in1                => s_in1(32,18),
			in2                => s_in2(32,18),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(18)
		);
	s_in1(32,18)            <= s_out1(33,18);
	s_in2(32,18)            <= s_out2(33,19);
	s_locks_lower_in(32,18) <= s_locks_lower_out(33,18);

		normal_cell_32_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,19),
			fetch              => s_fetch(32,19),
			data_in            => s_data_in(32,19),
			data_out           => s_data_out(32,19),
			out1               => s_out1(32,19),
			out2               => s_out2(32,19),
			lock_lower_row_out => s_locks_lower_out(32,19),
			lock_lower_row_in  => s_locks_lower_in(32,19),
			in1                => s_in1(32,19),
			in2                => s_in2(32,19),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(19)
		);
	s_in1(32,19)            <= s_out1(33,19);
	s_in2(32,19)            <= s_out2(33,20);
	s_locks_lower_in(32,19) <= s_locks_lower_out(33,19);

		normal_cell_32_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,20),
			fetch              => s_fetch(32,20),
			data_in            => s_data_in(32,20),
			data_out           => s_data_out(32,20),
			out1               => s_out1(32,20),
			out2               => s_out2(32,20),
			lock_lower_row_out => s_locks_lower_out(32,20),
			lock_lower_row_in  => s_locks_lower_in(32,20),
			in1                => s_in1(32,20),
			in2                => s_in2(32,20),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(20)
		);
	s_in1(32,20)            <= s_out1(33,20);
	s_in2(32,20)            <= s_out2(33,21);
	s_locks_lower_in(32,20) <= s_locks_lower_out(33,20);

		normal_cell_32_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,21),
			fetch              => s_fetch(32,21),
			data_in            => s_data_in(32,21),
			data_out           => s_data_out(32,21),
			out1               => s_out1(32,21),
			out2               => s_out2(32,21),
			lock_lower_row_out => s_locks_lower_out(32,21),
			lock_lower_row_in  => s_locks_lower_in(32,21),
			in1                => s_in1(32,21),
			in2                => s_in2(32,21),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(21)
		);
	s_in1(32,21)            <= s_out1(33,21);
	s_in2(32,21)            <= s_out2(33,22);
	s_locks_lower_in(32,21) <= s_locks_lower_out(33,21);

		normal_cell_32_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,22),
			fetch              => s_fetch(32,22),
			data_in            => s_data_in(32,22),
			data_out           => s_data_out(32,22),
			out1               => s_out1(32,22),
			out2               => s_out2(32,22),
			lock_lower_row_out => s_locks_lower_out(32,22),
			lock_lower_row_in  => s_locks_lower_in(32,22),
			in1                => s_in1(32,22),
			in2                => s_in2(32,22),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(22)
		);
	s_in1(32,22)            <= s_out1(33,22);
	s_in2(32,22)            <= s_out2(33,23);
	s_locks_lower_in(32,22) <= s_locks_lower_out(33,22);

		normal_cell_32_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,23),
			fetch              => s_fetch(32,23),
			data_in            => s_data_in(32,23),
			data_out           => s_data_out(32,23),
			out1               => s_out1(32,23),
			out2               => s_out2(32,23),
			lock_lower_row_out => s_locks_lower_out(32,23),
			lock_lower_row_in  => s_locks_lower_in(32,23),
			in1                => s_in1(32,23),
			in2                => s_in2(32,23),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(23)
		);
	s_in1(32,23)            <= s_out1(33,23);
	s_in2(32,23)            <= s_out2(33,24);
	s_locks_lower_in(32,23) <= s_locks_lower_out(33,23);

		normal_cell_32_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,24),
			fetch              => s_fetch(32,24),
			data_in            => s_data_in(32,24),
			data_out           => s_data_out(32,24),
			out1               => s_out1(32,24),
			out2               => s_out2(32,24),
			lock_lower_row_out => s_locks_lower_out(32,24),
			lock_lower_row_in  => s_locks_lower_in(32,24),
			in1                => s_in1(32,24),
			in2                => s_in2(32,24),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(24)
		);
	s_in1(32,24)            <= s_out1(33,24);
	s_in2(32,24)            <= s_out2(33,25);
	s_locks_lower_in(32,24) <= s_locks_lower_out(33,24);

		normal_cell_32_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,25),
			fetch              => s_fetch(32,25),
			data_in            => s_data_in(32,25),
			data_out           => s_data_out(32,25),
			out1               => s_out1(32,25),
			out2               => s_out2(32,25),
			lock_lower_row_out => s_locks_lower_out(32,25),
			lock_lower_row_in  => s_locks_lower_in(32,25),
			in1                => s_in1(32,25),
			in2                => s_in2(32,25),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(25)
		);
	s_in1(32,25)            <= s_out1(33,25);
	s_in2(32,25)            <= s_out2(33,26);
	s_locks_lower_in(32,25) <= s_locks_lower_out(33,25);

		normal_cell_32_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,26),
			fetch              => s_fetch(32,26),
			data_in            => s_data_in(32,26),
			data_out           => s_data_out(32,26),
			out1               => s_out1(32,26),
			out2               => s_out2(32,26),
			lock_lower_row_out => s_locks_lower_out(32,26),
			lock_lower_row_in  => s_locks_lower_in(32,26),
			in1                => s_in1(32,26),
			in2                => s_in2(32,26),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(26)
		);
	s_in1(32,26)            <= s_out1(33,26);
	s_in2(32,26)            <= s_out2(33,27);
	s_locks_lower_in(32,26) <= s_locks_lower_out(33,26);

		normal_cell_32_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,27),
			fetch              => s_fetch(32,27),
			data_in            => s_data_in(32,27),
			data_out           => s_data_out(32,27),
			out1               => s_out1(32,27),
			out2               => s_out2(32,27),
			lock_lower_row_out => s_locks_lower_out(32,27),
			lock_lower_row_in  => s_locks_lower_in(32,27),
			in1                => s_in1(32,27),
			in2                => s_in2(32,27),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(27)
		);
	s_in1(32,27)            <= s_out1(33,27);
	s_in2(32,27)            <= s_out2(33,28);
	s_locks_lower_in(32,27) <= s_locks_lower_out(33,27);

		normal_cell_32_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,28),
			fetch              => s_fetch(32,28),
			data_in            => s_data_in(32,28),
			data_out           => s_data_out(32,28),
			out1               => s_out1(32,28),
			out2               => s_out2(32,28),
			lock_lower_row_out => s_locks_lower_out(32,28),
			lock_lower_row_in  => s_locks_lower_in(32,28),
			in1                => s_in1(32,28),
			in2                => s_in2(32,28),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(28)
		);
	s_in1(32,28)            <= s_out1(33,28);
	s_in2(32,28)            <= s_out2(33,29);
	s_locks_lower_in(32,28) <= s_locks_lower_out(33,28);

		normal_cell_32_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,29),
			fetch              => s_fetch(32,29),
			data_in            => s_data_in(32,29),
			data_out           => s_data_out(32,29),
			out1               => s_out1(32,29),
			out2               => s_out2(32,29),
			lock_lower_row_out => s_locks_lower_out(32,29),
			lock_lower_row_in  => s_locks_lower_in(32,29),
			in1                => s_in1(32,29),
			in2                => s_in2(32,29),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(29)
		);
	s_in1(32,29)            <= s_out1(33,29);
	s_in2(32,29)            <= s_out2(33,30);
	s_locks_lower_in(32,29) <= s_locks_lower_out(33,29);

		normal_cell_32_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,30),
			fetch              => s_fetch(32,30),
			data_in            => s_data_in(32,30),
			data_out           => s_data_out(32,30),
			out1               => s_out1(32,30),
			out2               => s_out2(32,30),
			lock_lower_row_out => s_locks_lower_out(32,30),
			lock_lower_row_in  => s_locks_lower_in(32,30),
			in1                => s_in1(32,30),
			in2                => s_in2(32,30),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(30)
		);
	s_in1(32,30)            <= s_out1(33,30);
	s_in2(32,30)            <= s_out2(33,31);
	s_locks_lower_in(32,30) <= s_locks_lower_out(33,30);

		normal_cell_32_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,31),
			fetch              => s_fetch(32,31),
			data_in            => s_data_in(32,31),
			data_out           => s_data_out(32,31),
			out1               => s_out1(32,31),
			out2               => s_out2(32,31),
			lock_lower_row_out => s_locks_lower_out(32,31),
			lock_lower_row_in  => s_locks_lower_in(32,31),
			in1                => s_in1(32,31),
			in2                => s_in2(32,31),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(31)
		);
	s_in1(32,31)            <= s_out1(33,31);
	s_in2(32,31)            <= s_out2(33,32);
	s_locks_lower_in(32,31) <= s_locks_lower_out(33,31);

		normal_cell_32_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,32),
			fetch              => s_fetch(32,32),
			data_in            => s_data_in(32,32),
			data_out           => s_data_out(32,32),
			out1               => s_out1(32,32),
			out2               => s_out2(32,32),
			lock_lower_row_out => s_locks_lower_out(32,32),
			lock_lower_row_in  => s_locks_lower_in(32,32),
			in1                => s_in1(32,32),
			in2                => s_in2(32,32),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(32)
		);
	s_in1(32,32)            <= s_out1(33,32);
	s_in2(32,32)            <= s_out2(33,33);
	s_locks_lower_in(32,32) <= s_locks_lower_out(33,32);

		normal_cell_32_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,33),
			fetch              => s_fetch(32,33),
			data_in            => s_data_in(32,33),
			data_out           => s_data_out(32,33),
			out1               => s_out1(32,33),
			out2               => s_out2(32,33),
			lock_lower_row_out => s_locks_lower_out(32,33),
			lock_lower_row_in  => s_locks_lower_in(32,33),
			in1                => s_in1(32,33),
			in2                => s_in2(32,33),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(33)
		);
	s_in1(32,33)            <= s_out1(33,33);
	s_in2(32,33)            <= s_out2(33,34);
	s_locks_lower_in(32,33) <= s_locks_lower_out(33,33);

		normal_cell_32_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,34),
			fetch              => s_fetch(32,34),
			data_in            => s_data_in(32,34),
			data_out           => s_data_out(32,34),
			out1               => s_out1(32,34),
			out2               => s_out2(32,34),
			lock_lower_row_out => s_locks_lower_out(32,34),
			lock_lower_row_in  => s_locks_lower_in(32,34),
			in1                => s_in1(32,34),
			in2                => s_in2(32,34),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(34)
		);
	s_in1(32,34)            <= s_out1(33,34);
	s_in2(32,34)            <= s_out2(33,35);
	s_locks_lower_in(32,34) <= s_locks_lower_out(33,34);

		normal_cell_32_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,35),
			fetch              => s_fetch(32,35),
			data_in            => s_data_in(32,35),
			data_out           => s_data_out(32,35),
			out1               => s_out1(32,35),
			out2               => s_out2(32,35),
			lock_lower_row_out => s_locks_lower_out(32,35),
			lock_lower_row_in  => s_locks_lower_in(32,35),
			in1                => s_in1(32,35),
			in2                => s_in2(32,35),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(35)
		);
	s_in1(32,35)            <= s_out1(33,35);
	s_in2(32,35)            <= s_out2(33,36);
	s_locks_lower_in(32,35) <= s_locks_lower_out(33,35);

		normal_cell_32_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,36),
			fetch              => s_fetch(32,36),
			data_in            => s_data_in(32,36),
			data_out           => s_data_out(32,36),
			out1               => s_out1(32,36),
			out2               => s_out2(32,36),
			lock_lower_row_out => s_locks_lower_out(32,36),
			lock_lower_row_in  => s_locks_lower_in(32,36),
			in1                => s_in1(32,36),
			in2                => s_in2(32,36),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(36)
		);
	s_in1(32,36)            <= s_out1(33,36);
	s_in2(32,36)            <= s_out2(33,37);
	s_locks_lower_in(32,36) <= s_locks_lower_out(33,36);

		normal_cell_32_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,37),
			fetch              => s_fetch(32,37),
			data_in            => s_data_in(32,37),
			data_out           => s_data_out(32,37),
			out1               => s_out1(32,37),
			out2               => s_out2(32,37),
			lock_lower_row_out => s_locks_lower_out(32,37),
			lock_lower_row_in  => s_locks_lower_in(32,37),
			in1                => s_in1(32,37),
			in2                => s_in2(32,37),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(37)
		);
	s_in1(32,37)            <= s_out1(33,37);
	s_in2(32,37)            <= s_out2(33,38);
	s_locks_lower_in(32,37) <= s_locks_lower_out(33,37);

		normal_cell_32_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,38),
			fetch              => s_fetch(32,38),
			data_in            => s_data_in(32,38),
			data_out           => s_data_out(32,38),
			out1               => s_out1(32,38),
			out2               => s_out2(32,38),
			lock_lower_row_out => s_locks_lower_out(32,38),
			lock_lower_row_in  => s_locks_lower_in(32,38),
			in1                => s_in1(32,38),
			in2                => s_in2(32,38),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(38)
		);
	s_in1(32,38)            <= s_out1(33,38);
	s_in2(32,38)            <= s_out2(33,39);
	s_locks_lower_in(32,38) <= s_locks_lower_out(33,38);

		normal_cell_32_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,39),
			fetch              => s_fetch(32,39),
			data_in            => s_data_in(32,39),
			data_out           => s_data_out(32,39),
			out1               => s_out1(32,39),
			out2               => s_out2(32,39),
			lock_lower_row_out => s_locks_lower_out(32,39),
			lock_lower_row_in  => s_locks_lower_in(32,39),
			in1                => s_in1(32,39),
			in2                => s_in2(32,39),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(39)
		);
	s_in1(32,39)            <= s_out1(33,39);
	s_in2(32,39)            <= s_out2(33,40);
	s_locks_lower_in(32,39) <= s_locks_lower_out(33,39);

		normal_cell_32_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,40),
			fetch              => s_fetch(32,40),
			data_in            => s_data_in(32,40),
			data_out           => s_data_out(32,40),
			out1               => s_out1(32,40),
			out2               => s_out2(32,40),
			lock_lower_row_out => s_locks_lower_out(32,40),
			lock_lower_row_in  => s_locks_lower_in(32,40),
			in1                => s_in1(32,40),
			in2                => s_in2(32,40),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(40)
		);
	s_in1(32,40)            <= s_out1(33,40);
	s_in2(32,40)            <= s_out2(33,41);
	s_locks_lower_in(32,40) <= s_locks_lower_out(33,40);

		normal_cell_32_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,41),
			fetch              => s_fetch(32,41),
			data_in            => s_data_in(32,41),
			data_out           => s_data_out(32,41),
			out1               => s_out1(32,41),
			out2               => s_out2(32,41),
			lock_lower_row_out => s_locks_lower_out(32,41),
			lock_lower_row_in  => s_locks_lower_in(32,41),
			in1                => s_in1(32,41),
			in2                => s_in2(32,41),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(41)
		);
	s_in1(32,41)            <= s_out1(33,41);
	s_in2(32,41)            <= s_out2(33,42);
	s_locks_lower_in(32,41) <= s_locks_lower_out(33,41);

		normal_cell_32_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,42),
			fetch              => s_fetch(32,42),
			data_in            => s_data_in(32,42),
			data_out           => s_data_out(32,42),
			out1               => s_out1(32,42),
			out2               => s_out2(32,42),
			lock_lower_row_out => s_locks_lower_out(32,42),
			lock_lower_row_in  => s_locks_lower_in(32,42),
			in1                => s_in1(32,42),
			in2                => s_in2(32,42),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(42)
		);
	s_in1(32,42)            <= s_out1(33,42);
	s_in2(32,42)            <= s_out2(33,43);
	s_locks_lower_in(32,42) <= s_locks_lower_out(33,42);

		normal_cell_32_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,43),
			fetch              => s_fetch(32,43),
			data_in            => s_data_in(32,43),
			data_out           => s_data_out(32,43),
			out1               => s_out1(32,43),
			out2               => s_out2(32,43),
			lock_lower_row_out => s_locks_lower_out(32,43),
			lock_lower_row_in  => s_locks_lower_in(32,43),
			in1                => s_in1(32,43),
			in2                => s_in2(32,43),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(43)
		);
	s_in1(32,43)            <= s_out1(33,43);
	s_in2(32,43)            <= s_out2(33,44);
	s_locks_lower_in(32,43) <= s_locks_lower_out(33,43);

		normal_cell_32_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,44),
			fetch              => s_fetch(32,44),
			data_in            => s_data_in(32,44),
			data_out           => s_data_out(32,44),
			out1               => s_out1(32,44),
			out2               => s_out2(32,44),
			lock_lower_row_out => s_locks_lower_out(32,44),
			lock_lower_row_in  => s_locks_lower_in(32,44),
			in1                => s_in1(32,44),
			in2                => s_in2(32,44),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(44)
		);
	s_in1(32,44)            <= s_out1(33,44);
	s_in2(32,44)            <= s_out2(33,45);
	s_locks_lower_in(32,44) <= s_locks_lower_out(33,44);

		normal_cell_32_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,45),
			fetch              => s_fetch(32,45),
			data_in            => s_data_in(32,45),
			data_out           => s_data_out(32,45),
			out1               => s_out1(32,45),
			out2               => s_out2(32,45),
			lock_lower_row_out => s_locks_lower_out(32,45),
			lock_lower_row_in  => s_locks_lower_in(32,45),
			in1                => s_in1(32,45),
			in2                => s_in2(32,45),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(45)
		);
	s_in1(32,45)            <= s_out1(33,45);
	s_in2(32,45)            <= s_out2(33,46);
	s_locks_lower_in(32,45) <= s_locks_lower_out(33,45);

		normal_cell_32_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,46),
			fetch              => s_fetch(32,46),
			data_in            => s_data_in(32,46),
			data_out           => s_data_out(32,46),
			out1               => s_out1(32,46),
			out2               => s_out2(32,46),
			lock_lower_row_out => s_locks_lower_out(32,46),
			lock_lower_row_in  => s_locks_lower_in(32,46),
			in1                => s_in1(32,46),
			in2                => s_in2(32,46),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(46)
		);
	s_in1(32,46)            <= s_out1(33,46);
	s_in2(32,46)            <= s_out2(33,47);
	s_locks_lower_in(32,46) <= s_locks_lower_out(33,46);

		normal_cell_32_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,47),
			fetch              => s_fetch(32,47),
			data_in            => s_data_in(32,47),
			data_out           => s_data_out(32,47),
			out1               => s_out1(32,47),
			out2               => s_out2(32,47),
			lock_lower_row_out => s_locks_lower_out(32,47),
			lock_lower_row_in  => s_locks_lower_in(32,47),
			in1                => s_in1(32,47),
			in2                => s_in2(32,47),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(47)
		);
	s_in1(32,47)            <= s_out1(33,47);
	s_in2(32,47)            <= s_out2(33,48);
	s_locks_lower_in(32,47) <= s_locks_lower_out(33,47);

		normal_cell_32_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,48),
			fetch              => s_fetch(32,48),
			data_in            => s_data_in(32,48),
			data_out           => s_data_out(32,48),
			out1               => s_out1(32,48),
			out2               => s_out2(32,48),
			lock_lower_row_out => s_locks_lower_out(32,48),
			lock_lower_row_in  => s_locks_lower_in(32,48),
			in1                => s_in1(32,48),
			in2                => s_in2(32,48),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(48)
		);
	s_in1(32,48)            <= s_out1(33,48);
	s_in2(32,48)            <= s_out2(33,49);
	s_locks_lower_in(32,48) <= s_locks_lower_out(33,48);

		normal_cell_32_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,49),
			fetch              => s_fetch(32,49),
			data_in            => s_data_in(32,49),
			data_out           => s_data_out(32,49),
			out1               => s_out1(32,49),
			out2               => s_out2(32,49),
			lock_lower_row_out => s_locks_lower_out(32,49),
			lock_lower_row_in  => s_locks_lower_in(32,49),
			in1                => s_in1(32,49),
			in2                => s_in2(32,49),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(49)
		);
	s_in1(32,49)            <= s_out1(33,49);
	s_in2(32,49)            <= s_out2(33,50);
	s_locks_lower_in(32,49) <= s_locks_lower_out(33,49);

		normal_cell_32_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,50),
			fetch              => s_fetch(32,50),
			data_in            => s_data_in(32,50),
			data_out           => s_data_out(32,50),
			out1               => s_out1(32,50),
			out2               => s_out2(32,50),
			lock_lower_row_out => s_locks_lower_out(32,50),
			lock_lower_row_in  => s_locks_lower_in(32,50),
			in1                => s_in1(32,50),
			in2                => s_in2(32,50),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(50)
		);
	s_in1(32,50)            <= s_out1(33,50);
	s_in2(32,50)            <= s_out2(33,51);
	s_locks_lower_in(32,50) <= s_locks_lower_out(33,50);

		normal_cell_32_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,51),
			fetch              => s_fetch(32,51),
			data_in            => s_data_in(32,51),
			data_out           => s_data_out(32,51),
			out1               => s_out1(32,51),
			out2               => s_out2(32,51),
			lock_lower_row_out => s_locks_lower_out(32,51),
			lock_lower_row_in  => s_locks_lower_in(32,51),
			in1                => s_in1(32,51),
			in2                => s_in2(32,51),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(51)
		);
	s_in1(32,51)            <= s_out1(33,51);
	s_in2(32,51)            <= s_out2(33,52);
	s_locks_lower_in(32,51) <= s_locks_lower_out(33,51);

		normal_cell_32_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,52),
			fetch              => s_fetch(32,52),
			data_in            => s_data_in(32,52),
			data_out           => s_data_out(32,52),
			out1               => s_out1(32,52),
			out2               => s_out2(32,52),
			lock_lower_row_out => s_locks_lower_out(32,52),
			lock_lower_row_in  => s_locks_lower_in(32,52),
			in1                => s_in1(32,52),
			in2                => s_in2(32,52),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(52)
		);
	s_in1(32,52)            <= s_out1(33,52);
	s_in2(32,52)            <= s_out2(33,53);
	s_locks_lower_in(32,52) <= s_locks_lower_out(33,52);

		normal_cell_32_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,53),
			fetch              => s_fetch(32,53),
			data_in            => s_data_in(32,53),
			data_out           => s_data_out(32,53),
			out1               => s_out1(32,53),
			out2               => s_out2(32,53),
			lock_lower_row_out => s_locks_lower_out(32,53),
			lock_lower_row_in  => s_locks_lower_in(32,53),
			in1                => s_in1(32,53),
			in2                => s_in2(32,53),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(53)
		);
	s_in1(32,53)            <= s_out1(33,53);
	s_in2(32,53)            <= s_out2(33,54);
	s_locks_lower_in(32,53) <= s_locks_lower_out(33,53);

		normal_cell_32_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,54),
			fetch              => s_fetch(32,54),
			data_in            => s_data_in(32,54),
			data_out           => s_data_out(32,54),
			out1               => s_out1(32,54),
			out2               => s_out2(32,54),
			lock_lower_row_out => s_locks_lower_out(32,54),
			lock_lower_row_in  => s_locks_lower_in(32,54),
			in1                => s_in1(32,54),
			in2                => s_in2(32,54),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(54)
		);
	s_in1(32,54)            <= s_out1(33,54);
	s_in2(32,54)            <= s_out2(33,55);
	s_locks_lower_in(32,54) <= s_locks_lower_out(33,54);

		normal_cell_32_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,55),
			fetch              => s_fetch(32,55),
			data_in            => s_data_in(32,55),
			data_out           => s_data_out(32,55),
			out1               => s_out1(32,55),
			out2               => s_out2(32,55),
			lock_lower_row_out => s_locks_lower_out(32,55),
			lock_lower_row_in  => s_locks_lower_in(32,55),
			in1                => s_in1(32,55),
			in2                => s_in2(32,55),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(55)
		);
	s_in1(32,55)            <= s_out1(33,55);
	s_in2(32,55)            <= s_out2(33,56);
	s_locks_lower_in(32,55) <= s_locks_lower_out(33,55);

		normal_cell_32_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,56),
			fetch              => s_fetch(32,56),
			data_in            => s_data_in(32,56),
			data_out           => s_data_out(32,56),
			out1               => s_out1(32,56),
			out2               => s_out2(32,56),
			lock_lower_row_out => s_locks_lower_out(32,56),
			lock_lower_row_in  => s_locks_lower_in(32,56),
			in1                => s_in1(32,56),
			in2                => s_in2(32,56),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(56)
		);
	s_in1(32,56)            <= s_out1(33,56);
	s_in2(32,56)            <= s_out2(33,57);
	s_locks_lower_in(32,56) <= s_locks_lower_out(33,56);

		normal_cell_32_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,57),
			fetch              => s_fetch(32,57),
			data_in            => s_data_in(32,57),
			data_out           => s_data_out(32,57),
			out1               => s_out1(32,57),
			out2               => s_out2(32,57),
			lock_lower_row_out => s_locks_lower_out(32,57),
			lock_lower_row_in  => s_locks_lower_in(32,57),
			in1                => s_in1(32,57),
			in2                => s_in2(32,57),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(57)
		);
	s_in1(32,57)            <= s_out1(33,57);
	s_in2(32,57)            <= s_out2(33,58);
	s_locks_lower_in(32,57) <= s_locks_lower_out(33,57);

		normal_cell_32_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,58),
			fetch              => s_fetch(32,58),
			data_in            => s_data_in(32,58),
			data_out           => s_data_out(32,58),
			out1               => s_out1(32,58),
			out2               => s_out2(32,58),
			lock_lower_row_out => s_locks_lower_out(32,58),
			lock_lower_row_in  => s_locks_lower_in(32,58),
			in1                => s_in1(32,58),
			in2                => s_in2(32,58),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(58)
		);
	s_in1(32,58)            <= s_out1(33,58);
	s_in2(32,58)            <= s_out2(33,59);
	s_locks_lower_in(32,58) <= s_locks_lower_out(33,58);

		normal_cell_32_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,59),
			fetch              => s_fetch(32,59),
			data_in            => s_data_in(32,59),
			data_out           => s_data_out(32,59),
			out1               => s_out1(32,59),
			out2               => s_out2(32,59),
			lock_lower_row_out => s_locks_lower_out(32,59),
			lock_lower_row_in  => s_locks_lower_in(32,59),
			in1                => s_in1(32,59),
			in2                => s_in2(32,59),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(59)
		);
	s_in1(32,59)            <= s_out1(33,59);
	s_in2(32,59)            <= s_out2(33,60);
	s_locks_lower_in(32,59) <= s_locks_lower_out(33,59);

		last_col_cell_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(32,60),
			fetch              => s_fetch(32,60),
			data_in            => s_data_in(32,60),
			data_out           => s_data_out(32,60),
			out1               => s_out1(32,60),
			out2               => s_out2(32,60),
			lock_lower_row_out => s_locks_lower_out(32,60),
			lock_lower_row_in  => s_locks_lower_in(32,60),
			in1                => s_in1(32,60),
			in2                => (others => '0'),
			lock_row           => s_locks(32),
			piv_found          => s_piv_found,
			row_data           => s_row_data(32),
			col_data           => s_col_data(60)
		);
	s_in1(32,60)            <= s_out1(33,60);
	s_locks_lower_in(32,60) <= s_locks_lower_out(33,60);

		normal_cell_33_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,1),
			fetch              => s_fetch(33,1),
			data_in            => s_data_in(33,1),
			data_out           => s_data_out(33,1),
			out1               => s_out1(33,1),
			out2               => s_out2(33,1),
			lock_lower_row_out => s_locks_lower_out(33,1),
			lock_lower_row_in  => s_locks_lower_in(33,1),
			in1                => s_in1(33,1),
			in2                => s_in2(33,1),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(1)
		);
	s_in1(33,1)            <= s_out1(34,1);
	s_in2(33,1)            <= s_out2(34,2);
	s_locks_lower_in(33,1) <= s_locks_lower_out(34,1);

		normal_cell_33_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,2),
			fetch              => s_fetch(33,2),
			data_in            => s_data_in(33,2),
			data_out           => s_data_out(33,2),
			out1               => s_out1(33,2),
			out2               => s_out2(33,2),
			lock_lower_row_out => s_locks_lower_out(33,2),
			lock_lower_row_in  => s_locks_lower_in(33,2),
			in1                => s_in1(33,2),
			in2                => s_in2(33,2),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(2)
		);
	s_in1(33,2)            <= s_out1(34,2);
	s_in2(33,2)            <= s_out2(34,3);
	s_locks_lower_in(33,2) <= s_locks_lower_out(34,2);

		normal_cell_33_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,3),
			fetch              => s_fetch(33,3),
			data_in            => s_data_in(33,3),
			data_out           => s_data_out(33,3),
			out1               => s_out1(33,3),
			out2               => s_out2(33,3),
			lock_lower_row_out => s_locks_lower_out(33,3),
			lock_lower_row_in  => s_locks_lower_in(33,3),
			in1                => s_in1(33,3),
			in2                => s_in2(33,3),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(3)
		);
	s_in1(33,3)            <= s_out1(34,3);
	s_in2(33,3)            <= s_out2(34,4);
	s_locks_lower_in(33,3) <= s_locks_lower_out(34,3);

		normal_cell_33_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,4),
			fetch              => s_fetch(33,4),
			data_in            => s_data_in(33,4),
			data_out           => s_data_out(33,4),
			out1               => s_out1(33,4),
			out2               => s_out2(33,4),
			lock_lower_row_out => s_locks_lower_out(33,4),
			lock_lower_row_in  => s_locks_lower_in(33,4),
			in1                => s_in1(33,4),
			in2                => s_in2(33,4),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(4)
		);
	s_in1(33,4)            <= s_out1(34,4);
	s_in2(33,4)            <= s_out2(34,5);
	s_locks_lower_in(33,4) <= s_locks_lower_out(34,4);

		normal_cell_33_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,5),
			fetch              => s_fetch(33,5),
			data_in            => s_data_in(33,5),
			data_out           => s_data_out(33,5),
			out1               => s_out1(33,5),
			out2               => s_out2(33,5),
			lock_lower_row_out => s_locks_lower_out(33,5),
			lock_lower_row_in  => s_locks_lower_in(33,5),
			in1                => s_in1(33,5),
			in2                => s_in2(33,5),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(5)
		);
	s_in1(33,5)            <= s_out1(34,5);
	s_in2(33,5)            <= s_out2(34,6);
	s_locks_lower_in(33,5) <= s_locks_lower_out(34,5);

		normal_cell_33_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,6),
			fetch              => s_fetch(33,6),
			data_in            => s_data_in(33,6),
			data_out           => s_data_out(33,6),
			out1               => s_out1(33,6),
			out2               => s_out2(33,6),
			lock_lower_row_out => s_locks_lower_out(33,6),
			lock_lower_row_in  => s_locks_lower_in(33,6),
			in1                => s_in1(33,6),
			in2                => s_in2(33,6),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(6)
		);
	s_in1(33,6)            <= s_out1(34,6);
	s_in2(33,6)            <= s_out2(34,7);
	s_locks_lower_in(33,6) <= s_locks_lower_out(34,6);

		normal_cell_33_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,7),
			fetch              => s_fetch(33,7),
			data_in            => s_data_in(33,7),
			data_out           => s_data_out(33,7),
			out1               => s_out1(33,7),
			out2               => s_out2(33,7),
			lock_lower_row_out => s_locks_lower_out(33,7),
			lock_lower_row_in  => s_locks_lower_in(33,7),
			in1                => s_in1(33,7),
			in2                => s_in2(33,7),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(7)
		);
	s_in1(33,7)            <= s_out1(34,7);
	s_in2(33,7)            <= s_out2(34,8);
	s_locks_lower_in(33,7) <= s_locks_lower_out(34,7);

		normal_cell_33_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,8),
			fetch              => s_fetch(33,8),
			data_in            => s_data_in(33,8),
			data_out           => s_data_out(33,8),
			out1               => s_out1(33,8),
			out2               => s_out2(33,8),
			lock_lower_row_out => s_locks_lower_out(33,8),
			lock_lower_row_in  => s_locks_lower_in(33,8),
			in1                => s_in1(33,8),
			in2                => s_in2(33,8),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(8)
		);
	s_in1(33,8)            <= s_out1(34,8);
	s_in2(33,8)            <= s_out2(34,9);
	s_locks_lower_in(33,8) <= s_locks_lower_out(34,8);

		normal_cell_33_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,9),
			fetch              => s_fetch(33,9),
			data_in            => s_data_in(33,9),
			data_out           => s_data_out(33,9),
			out1               => s_out1(33,9),
			out2               => s_out2(33,9),
			lock_lower_row_out => s_locks_lower_out(33,9),
			lock_lower_row_in  => s_locks_lower_in(33,9),
			in1                => s_in1(33,9),
			in2                => s_in2(33,9),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(9)
		);
	s_in1(33,9)            <= s_out1(34,9);
	s_in2(33,9)            <= s_out2(34,10);
	s_locks_lower_in(33,9) <= s_locks_lower_out(34,9);

		normal_cell_33_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,10),
			fetch              => s_fetch(33,10),
			data_in            => s_data_in(33,10),
			data_out           => s_data_out(33,10),
			out1               => s_out1(33,10),
			out2               => s_out2(33,10),
			lock_lower_row_out => s_locks_lower_out(33,10),
			lock_lower_row_in  => s_locks_lower_in(33,10),
			in1                => s_in1(33,10),
			in2                => s_in2(33,10),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(10)
		);
	s_in1(33,10)            <= s_out1(34,10);
	s_in2(33,10)            <= s_out2(34,11);
	s_locks_lower_in(33,10) <= s_locks_lower_out(34,10);

		normal_cell_33_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,11),
			fetch              => s_fetch(33,11),
			data_in            => s_data_in(33,11),
			data_out           => s_data_out(33,11),
			out1               => s_out1(33,11),
			out2               => s_out2(33,11),
			lock_lower_row_out => s_locks_lower_out(33,11),
			lock_lower_row_in  => s_locks_lower_in(33,11),
			in1                => s_in1(33,11),
			in2                => s_in2(33,11),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(11)
		);
	s_in1(33,11)            <= s_out1(34,11);
	s_in2(33,11)            <= s_out2(34,12);
	s_locks_lower_in(33,11) <= s_locks_lower_out(34,11);

		normal_cell_33_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,12),
			fetch              => s_fetch(33,12),
			data_in            => s_data_in(33,12),
			data_out           => s_data_out(33,12),
			out1               => s_out1(33,12),
			out2               => s_out2(33,12),
			lock_lower_row_out => s_locks_lower_out(33,12),
			lock_lower_row_in  => s_locks_lower_in(33,12),
			in1                => s_in1(33,12),
			in2                => s_in2(33,12),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(12)
		);
	s_in1(33,12)            <= s_out1(34,12);
	s_in2(33,12)            <= s_out2(34,13);
	s_locks_lower_in(33,12) <= s_locks_lower_out(34,12);

		normal_cell_33_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,13),
			fetch              => s_fetch(33,13),
			data_in            => s_data_in(33,13),
			data_out           => s_data_out(33,13),
			out1               => s_out1(33,13),
			out2               => s_out2(33,13),
			lock_lower_row_out => s_locks_lower_out(33,13),
			lock_lower_row_in  => s_locks_lower_in(33,13),
			in1                => s_in1(33,13),
			in2                => s_in2(33,13),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(13)
		);
	s_in1(33,13)            <= s_out1(34,13);
	s_in2(33,13)            <= s_out2(34,14);
	s_locks_lower_in(33,13) <= s_locks_lower_out(34,13);

		normal_cell_33_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,14),
			fetch              => s_fetch(33,14),
			data_in            => s_data_in(33,14),
			data_out           => s_data_out(33,14),
			out1               => s_out1(33,14),
			out2               => s_out2(33,14),
			lock_lower_row_out => s_locks_lower_out(33,14),
			lock_lower_row_in  => s_locks_lower_in(33,14),
			in1                => s_in1(33,14),
			in2                => s_in2(33,14),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(14)
		);
	s_in1(33,14)            <= s_out1(34,14);
	s_in2(33,14)            <= s_out2(34,15);
	s_locks_lower_in(33,14) <= s_locks_lower_out(34,14);

		normal_cell_33_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,15),
			fetch              => s_fetch(33,15),
			data_in            => s_data_in(33,15),
			data_out           => s_data_out(33,15),
			out1               => s_out1(33,15),
			out2               => s_out2(33,15),
			lock_lower_row_out => s_locks_lower_out(33,15),
			lock_lower_row_in  => s_locks_lower_in(33,15),
			in1                => s_in1(33,15),
			in2                => s_in2(33,15),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(15)
		);
	s_in1(33,15)            <= s_out1(34,15);
	s_in2(33,15)            <= s_out2(34,16);
	s_locks_lower_in(33,15) <= s_locks_lower_out(34,15);

		normal_cell_33_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,16),
			fetch              => s_fetch(33,16),
			data_in            => s_data_in(33,16),
			data_out           => s_data_out(33,16),
			out1               => s_out1(33,16),
			out2               => s_out2(33,16),
			lock_lower_row_out => s_locks_lower_out(33,16),
			lock_lower_row_in  => s_locks_lower_in(33,16),
			in1                => s_in1(33,16),
			in2                => s_in2(33,16),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(16)
		);
	s_in1(33,16)            <= s_out1(34,16);
	s_in2(33,16)            <= s_out2(34,17);
	s_locks_lower_in(33,16) <= s_locks_lower_out(34,16);

		normal_cell_33_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,17),
			fetch              => s_fetch(33,17),
			data_in            => s_data_in(33,17),
			data_out           => s_data_out(33,17),
			out1               => s_out1(33,17),
			out2               => s_out2(33,17),
			lock_lower_row_out => s_locks_lower_out(33,17),
			lock_lower_row_in  => s_locks_lower_in(33,17),
			in1                => s_in1(33,17),
			in2                => s_in2(33,17),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(17)
		);
	s_in1(33,17)            <= s_out1(34,17);
	s_in2(33,17)            <= s_out2(34,18);
	s_locks_lower_in(33,17) <= s_locks_lower_out(34,17);

		normal_cell_33_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,18),
			fetch              => s_fetch(33,18),
			data_in            => s_data_in(33,18),
			data_out           => s_data_out(33,18),
			out1               => s_out1(33,18),
			out2               => s_out2(33,18),
			lock_lower_row_out => s_locks_lower_out(33,18),
			lock_lower_row_in  => s_locks_lower_in(33,18),
			in1                => s_in1(33,18),
			in2                => s_in2(33,18),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(18)
		);
	s_in1(33,18)            <= s_out1(34,18);
	s_in2(33,18)            <= s_out2(34,19);
	s_locks_lower_in(33,18) <= s_locks_lower_out(34,18);

		normal_cell_33_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,19),
			fetch              => s_fetch(33,19),
			data_in            => s_data_in(33,19),
			data_out           => s_data_out(33,19),
			out1               => s_out1(33,19),
			out2               => s_out2(33,19),
			lock_lower_row_out => s_locks_lower_out(33,19),
			lock_lower_row_in  => s_locks_lower_in(33,19),
			in1                => s_in1(33,19),
			in2                => s_in2(33,19),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(19)
		);
	s_in1(33,19)            <= s_out1(34,19);
	s_in2(33,19)            <= s_out2(34,20);
	s_locks_lower_in(33,19) <= s_locks_lower_out(34,19);

		normal_cell_33_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,20),
			fetch              => s_fetch(33,20),
			data_in            => s_data_in(33,20),
			data_out           => s_data_out(33,20),
			out1               => s_out1(33,20),
			out2               => s_out2(33,20),
			lock_lower_row_out => s_locks_lower_out(33,20),
			lock_lower_row_in  => s_locks_lower_in(33,20),
			in1                => s_in1(33,20),
			in2                => s_in2(33,20),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(20)
		);
	s_in1(33,20)            <= s_out1(34,20);
	s_in2(33,20)            <= s_out2(34,21);
	s_locks_lower_in(33,20) <= s_locks_lower_out(34,20);

		normal_cell_33_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,21),
			fetch              => s_fetch(33,21),
			data_in            => s_data_in(33,21),
			data_out           => s_data_out(33,21),
			out1               => s_out1(33,21),
			out2               => s_out2(33,21),
			lock_lower_row_out => s_locks_lower_out(33,21),
			lock_lower_row_in  => s_locks_lower_in(33,21),
			in1                => s_in1(33,21),
			in2                => s_in2(33,21),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(21)
		);
	s_in1(33,21)            <= s_out1(34,21);
	s_in2(33,21)            <= s_out2(34,22);
	s_locks_lower_in(33,21) <= s_locks_lower_out(34,21);

		normal_cell_33_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,22),
			fetch              => s_fetch(33,22),
			data_in            => s_data_in(33,22),
			data_out           => s_data_out(33,22),
			out1               => s_out1(33,22),
			out2               => s_out2(33,22),
			lock_lower_row_out => s_locks_lower_out(33,22),
			lock_lower_row_in  => s_locks_lower_in(33,22),
			in1                => s_in1(33,22),
			in2                => s_in2(33,22),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(22)
		);
	s_in1(33,22)            <= s_out1(34,22);
	s_in2(33,22)            <= s_out2(34,23);
	s_locks_lower_in(33,22) <= s_locks_lower_out(34,22);

		normal_cell_33_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,23),
			fetch              => s_fetch(33,23),
			data_in            => s_data_in(33,23),
			data_out           => s_data_out(33,23),
			out1               => s_out1(33,23),
			out2               => s_out2(33,23),
			lock_lower_row_out => s_locks_lower_out(33,23),
			lock_lower_row_in  => s_locks_lower_in(33,23),
			in1                => s_in1(33,23),
			in2                => s_in2(33,23),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(23)
		);
	s_in1(33,23)            <= s_out1(34,23);
	s_in2(33,23)            <= s_out2(34,24);
	s_locks_lower_in(33,23) <= s_locks_lower_out(34,23);

		normal_cell_33_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,24),
			fetch              => s_fetch(33,24),
			data_in            => s_data_in(33,24),
			data_out           => s_data_out(33,24),
			out1               => s_out1(33,24),
			out2               => s_out2(33,24),
			lock_lower_row_out => s_locks_lower_out(33,24),
			lock_lower_row_in  => s_locks_lower_in(33,24),
			in1                => s_in1(33,24),
			in2                => s_in2(33,24),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(24)
		);
	s_in1(33,24)            <= s_out1(34,24);
	s_in2(33,24)            <= s_out2(34,25);
	s_locks_lower_in(33,24) <= s_locks_lower_out(34,24);

		normal_cell_33_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,25),
			fetch              => s_fetch(33,25),
			data_in            => s_data_in(33,25),
			data_out           => s_data_out(33,25),
			out1               => s_out1(33,25),
			out2               => s_out2(33,25),
			lock_lower_row_out => s_locks_lower_out(33,25),
			lock_lower_row_in  => s_locks_lower_in(33,25),
			in1                => s_in1(33,25),
			in2                => s_in2(33,25),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(25)
		);
	s_in1(33,25)            <= s_out1(34,25);
	s_in2(33,25)            <= s_out2(34,26);
	s_locks_lower_in(33,25) <= s_locks_lower_out(34,25);

		normal_cell_33_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,26),
			fetch              => s_fetch(33,26),
			data_in            => s_data_in(33,26),
			data_out           => s_data_out(33,26),
			out1               => s_out1(33,26),
			out2               => s_out2(33,26),
			lock_lower_row_out => s_locks_lower_out(33,26),
			lock_lower_row_in  => s_locks_lower_in(33,26),
			in1                => s_in1(33,26),
			in2                => s_in2(33,26),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(26)
		);
	s_in1(33,26)            <= s_out1(34,26);
	s_in2(33,26)            <= s_out2(34,27);
	s_locks_lower_in(33,26) <= s_locks_lower_out(34,26);

		normal_cell_33_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,27),
			fetch              => s_fetch(33,27),
			data_in            => s_data_in(33,27),
			data_out           => s_data_out(33,27),
			out1               => s_out1(33,27),
			out2               => s_out2(33,27),
			lock_lower_row_out => s_locks_lower_out(33,27),
			lock_lower_row_in  => s_locks_lower_in(33,27),
			in1                => s_in1(33,27),
			in2                => s_in2(33,27),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(27)
		);
	s_in1(33,27)            <= s_out1(34,27);
	s_in2(33,27)            <= s_out2(34,28);
	s_locks_lower_in(33,27) <= s_locks_lower_out(34,27);

		normal_cell_33_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,28),
			fetch              => s_fetch(33,28),
			data_in            => s_data_in(33,28),
			data_out           => s_data_out(33,28),
			out1               => s_out1(33,28),
			out2               => s_out2(33,28),
			lock_lower_row_out => s_locks_lower_out(33,28),
			lock_lower_row_in  => s_locks_lower_in(33,28),
			in1                => s_in1(33,28),
			in2                => s_in2(33,28),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(28)
		);
	s_in1(33,28)            <= s_out1(34,28);
	s_in2(33,28)            <= s_out2(34,29);
	s_locks_lower_in(33,28) <= s_locks_lower_out(34,28);

		normal_cell_33_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,29),
			fetch              => s_fetch(33,29),
			data_in            => s_data_in(33,29),
			data_out           => s_data_out(33,29),
			out1               => s_out1(33,29),
			out2               => s_out2(33,29),
			lock_lower_row_out => s_locks_lower_out(33,29),
			lock_lower_row_in  => s_locks_lower_in(33,29),
			in1                => s_in1(33,29),
			in2                => s_in2(33,29),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(29)
		);
	s_in1(33,29)            <= s_out1(34,29);
	s_in2(33,29)            <= s_out2(34,30);
	s_locks_lower_in(33,29) <= s_locks_lower_out(34,29);

		normal_cell_33_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,30),
			fetch              => s_fetch(33,30),
			data_in            => s_data_in(33,30),
			data_out           => s_data_out(33,30),
			out1               => s_out1(33,30),
			out2               => s_out2(33,30),
			lock_lower_row_out => s_locks_lower_out(33,30),
			lock_lower_row_in  => s_locks_lower_in(33,30),
			in1                => s_in1(33,30),
			in2                => s_in2(33,30),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(30)
		);
	s_in1(33,30)            <= s_out1(34,30);
	s_in2(33,30)            <= s_out2(34,31);
	s_locks_lower_in(33,30) <= s_locks_lower_out(34,30);

		normal_cell_33_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,31),
			fetch              => s_fetch(33,31),
			data_in            => s_data_in(33,31),
			data_out           => s_data_out(33,31),
			out1               => s_out1(33,31),
			out2               => s_out2(33,31),
			lock_lower_row_out => s_locks_lower_out(33,31),
			lock_lower_row_in  => s_locks_lower_in(33,31),
			in1                => s_in1(33,31),
			in2                => s_in2(33,31),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(31)
		);
	s_in1(33,31)            <= s_out1(34,31);
	s_in2(33,31)            <= s_out2(34,32);
	s_locks_lower_in(33,31) <= s_locks_lower_out(34,31);

		normal_cell_33_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,32),
			fetch              => s_fetch(33,32),
			data_in            => s_data_in(33,32),
			data_out           => s_data_out(33,32),
			out1               => s_out1(33,32),
			out2               => s_out2(33,32),
			lock_lower_row_out => s_locks_lower_out(33,32),
			lock_lower_row_in  => s_locks_lower_in(33,32),
			in1                => s_in1(33,32),
			in2                => s_in2(33,32),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(32)
		);
	s_in1(33,32)            <= s_out1(34,32);
	s_in2(33,32)            <= s_out2(34,33);
	s_locks_lower_in(33,32) <= s_locks_lower_out(34,32);

		normal_cell_33_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,33),
			fetch              => s_fetch(33,33),
			data_in            => s_data_in(33,33),
			data_out           => s_data_out(33,33),
			out1               => s_out1(33,33),
			out2               => s_out2(33,33),
			lock_lower_row_out => s_locks_lower_out(33,33),
			lock_lower_row_in  => s_locks_lower_in(33,33),
			in1                => s_in1(33,33),
			in2                => s_in2(33,33),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(33)
		);
	s_in1(33,33)            <= s_out1(34,33);
	s_in2(33,33)            <= s_out2(34,34);
	s_locks_lower_in(33,33) <= s_locks_lower_out(34,33);

		normal_cell_33_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,34),
			fetch              => s_fetch(33,34),
			data_in            => s_data_in(33,34),
			data_out           => s_data_out(33,34),
			out1               => s_out1(33,34),
			out2               => s_out2(33,34),
			lock_lower_row_out => s_locks_lower_out(33,34),
			lock_lower_row_in  => s_locks_lower_in(33,34),
			in1                => s_in1(33,34),
			in2                => s_in2(33,34),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(34)
		);
	s_in1(33,34)            <= s_out1(34,34);
	s_in2(33,34)            <= s_out2(34,35);
	s_locks_lower_in(33,34) <= s_locks_lower_out(34,34);

		normal_cell_33_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,35),
			fetch              => s_fetch(33,35),
			data_in            => s_data_in(33,35),
			data_out           => s_data_out(33,35),
			out1               => s_out1(33,35),
			out2               => s_out2(33,35),
			lock_lower_row_out => s_locks_lower_out(33,35),
			lock_lower_row_in  => s_locks_lower_in(33,35),
			in1                => s_in1(33,35),
			in2                => s_in2(33,35),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(35)
		);
	s_in1(33,35)            <= s_out1(34,35);
	s_in2(33,35)            <= s_out2(34,36);
	s_locks_lower_in(33,35) <= s_locks_lower_out(34,35);

		normal_cell_33_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,36),
			fetch              => s_fetch(33,36),
			data_in            => s_data_in(33,36),
			data_out           => s_data_out(33,36),
			out1               => s_out1(33,36),
			out2               => s_out2(33,36),
			lock_lower_row_out => s_locks_lower_out(33,36),
			lock_lower_row_in  => s_locks_lower_in(33,36),
			in1                => s_in1(33,36),
			in2                => s_in2(33,36),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(36)
		);
	s_in1(33,36)            <= s_out1(34,36);
	s_in2(33,36)            <= s_out2(34,37);
	s_locks_lower_in(33,36) <= s_locks_lower_out(34,36);

		normal_cell_33_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,37),
			fetch              => s_fetch(33,37),
			data_in            => s_data_in(33,37),
			data_out           => s_data_out(33,37),
			out1               => s_out1(33,37),
			out2               => s_out2(33,37),
			lock_lower_row_out => s_locks_lower_out(33,37),
			lock_lower_row_in  => s_locks_lower_in(33,37),
			in1                => s_in1(33,37),
			in2                => s_in2(33,37),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(37)
		);
	s_in1(33,37)            <= s_out1(34,37);
	s_in2(33,37)            <= s_out2(34,38);
	s_locks_lower_in(33,37) <= s_locks_lower_out(34,37);

		normal_cell_33_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,38),
			fetch              => s_fetch(33,38),
			data_in            => s_data_in(33,38),
			data_out           => s_data_out(33,38),
			out1               => s_out1(33,38),
			out2               => s_out2(33,38),
			lock_lower_row_out => s_locks_lower_out(33,38),
			lock_lower_row_in  => s_locks_lower_in(33,38),
			in1                => s_in1(33,38),
			in2                => s_in2(33,38),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(38)
		);
	s_in1(33,38)            <= s_out1(34,38);
	s_in2(33,38)            <= s_out2(34,39);
	s_locks_lower_in(33,38) <= s_locks_lower_out(34,38);

		normal_cell_33_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,39),
			fetch              => s_fetch(33,39),
			data_in            => s_data_in(33,39),
			data_out           => s_data_out(33,39),
			out1               => s_out1(33,39),
			out2               => s_out2(33,39),
			lock_lower_row_out => s_locks_lower_out(33,39),
			lock_lower_row_in  => s_locks_lower_in(33,39),
			in1                => s_in1(33,39),
			in2                => s_in2(33,39),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(39)
		);
	s_in1(33,39)            <= s_out1(34,39);
	s_in2(33,39)            <= s_out2(34,40);
	s_locks_lower_in(33,39) <= s_locks_lower_out(34,39);

		normal_cell_33_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,40),
			fetch              => s_fetch(33,40),
			data_in            => s_data_in(33,40),
			data_out           => s_data_out(33,40),
			out1               => s_out1(33,40),
			out2               => s_out2(33,40),
			lock_lower_row_out => s_locks_lower_out(33,40),
			lock_lower_row_in  => s_locks_lower_in(33,40),
			in1                => s_in1(33,40),
			in2                => s_in2(33,40),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(40)
		);
	s_in1(33,40)            <= s_out1(34,40);
	s_in2(33,40)            <= s_out2(34,41);
	s_locks_lower_in(33,40) <= s_locks_lower_out(34,40);

		normal_cell_33_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,41),
			fetch              => s_fetch(33,41),
			data_in            => s_data_in(33,41),
			data_out           => s_data_out(33,41),
			out1               => s_out1(33,41),
			out2               => s_out2(33,41),
			lock_lower_row_out => s_locks_lower_out(33,41),
			lock_lower_row_in  => s_locks_lower_in(33,41),
			in1                => s_in1(33,41),
			in2                => s_in2(33,41),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(41)
		);
	s_in1(33,41)            <= s_out1(34,41);
	s_in2(33,41)            <= s_out2(34,42);
	s_locks_lower_in(33,41) <= s_locks_lower_out(34,41);

		normal_cell_33_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,42),
			fetch              => s_fetch(33,42),
			data_in            => s_data_in(33,42),
			data_out           => s_data_out(33,42),
			out1               => s_out1(33,42),
			out2               => s_out2(33,42),
			lock_lower_row_out => s_locks_lower_out(33,42),
			lock_lower_row_in  => s_locks_lower_in(33,42),
			in1                => s_in1(33,42),
			in2                => s_in2(33,42),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(42)
		);
	s_in1(33,42)            <= s_out1(34,42);
	s_in2(33,42)            <= s_out2(34,43);
	s_locks_lower_in(33,42) <= s_locks_lower_out(34,42);

		normal_cell_33_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,43),
			fetch              => s_fetch(33,43),
			data_in            => s_data_in(33,43),
			data_out           => s_data_out(33,43),
			out1               => s_out1(33,43),
			out2               => s_out2(33,43),
			lock_lower_row_out => s_locks_lower_out(33,43),
			lock_lower_row_in  => s_locks_lower_in(33,43),
			in1                => s_in1(33,43),
			in2                => s_in2(33,43),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(43)
		);
	s_in1(33,43)            <= s_out1(34,43);
	s_in2(33,43)            <= s_out2(34,44);
	s_locks_lower_in(33,43) <= s_locks_lower_out(34,43);

		normal_cell_33_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,44),
			fetch              => s_fetch(33,44),
			data_in            => s_data_in(33,44),
			data_out           => s_data_out(33,44),
			out1               => s_out1(33,44),
			out2               => s_out2(33,44),
			lock_lower_row_out => s_locks_lower_out(33,44),
			lock_lower_row_in  => s_locks_lower_in(33,44),
			in1                => s_in1(33,44),
			in2                => s_in2(33,44),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(44)
		);
	s_in1(33,44)            <= s_out1(34,44);
	s_in2(33,44)            <= s_out2(34,45);
	s_locks_lower_in(33,44) <= s_locks_lower_out(34,44);

		normal_cell_33_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,45),
			fetch              => s_fetch(33,45),
			data_in            => s_data_in(33,45),
			data_out           => s_data_out(33,45),
			out1               => s_out1(33,45),
			out2               => s_out2(33,45),
			lock_lower_row_out => s_locks_lower_out(33,45),
			lock_lower_row_in  => s_locks_lower_in(33,45),
			in1                => s_in1(33,45),
			in2                => s_in2(33,45),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(45)
		);
	s_in1(33,45)            <= s_out1(34,45);
	s_in2(33,45)            <= s_out2(34,46);
	s_locks_lower_in(33,45) <= s_locks_lower_out(34,45);

		normal_cell_33_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,46),
			fetch              => s_fetch(33,46),
			data_in            => s_data_in(33,46),
			data_out           => s_data_out(33,46),
			out1               => s_out1(33,46),
			out2               => s_out2(33,46),
			lock_lower_row_out => s_locks_lower_out(33,46),
			lock_lower_row_in  => s_locks_lower_in(33,46),
			in1                => s_in1(33,46),
			in2                => s_in2(33,46),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(46)
		);
	s_in1(33,46)            <= s_out1(34,46);
	s_in2(33,46)            <= s_out2(34,47);
	s_locks_lower_in(33,46) <= s_locks_lower_out(34,46);

		normal_cell_33_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,47),
			fetch              => s_fetch(33,47),
			data_in            => s_data_in(33,47),
			data_out           => s_data_out(33,47),
			out1               => s_out1(33,47),
			out2               => s_out2(33,47),
			lock_lower_row_out => s_locks_lower_out(33,47),
			lock_lower_row_in  => s_locks_lower_in(33,47),
			in1                => s_in1(33,47),
			in2                => s_in2(33,47),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(47)
		);
	s_in1(33,47)            <= s_out1(34,47);
	s_in2(33,47)            <= s_out2(34,48);
	s_locks_lower_in(33,47) <= s_locks_lower_out(34,47);

		normal_cell_33_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,48),
			fetch              => s_fetch(33,48),
			data_in            => s_data_in(33,48),
			data_out           => s_data_out(33,48),
			out1               => s_out1(33,48),
			out2               => s_out2(33,48),
			lock_lower_row_out => s_locks_lower_out(33,48),
			lock_lower_row_in  => s_locks_lower_in(33,48),
			in1                => s_in1(33,48),
			in2                => s_in2(33,48),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(48)
		);
	s_in1(33,48)            <= s_out1(34,48);
	s_in2(33,48)            <= s_out2(34,49);
	s_locks_lower_in(33,48) <= s_locks_lower_out(34,48);

		normal_cell_33_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,49),
			fetch              => s_fetch(33,49),
			data_in            => s_data_in(33,49),
			data_out           => s_data_out(33,49),
			out1               => s_out1(33,49),
			out2               => s_out2(33,49),
			lock_lower_row_out => s_locks_lower_out(33,49),
			lock_lower_row_in  => s_locks_lower_in(33,49),
			in1                => s_in1(33,49),
			in2                => s_in2(33,49),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(49)
		);
	s_in1(33,49)            <= s_out1(34,49);
	s_in2(33,49)            <= s_out2(34,50);
	s_locks_lower_in(33,49) <= s_locks_lower_out(34,49);

		normal_cell_33_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,50),
			fetch              => s_fetch(33,50),
			data_in            => s_data_in(33,50),
			data_out           => s_data_out(33,50),
			out1               => s_out1(33,50),
			out2               => s_out2(33,50),
			lock_lower_row_out => s_locks_lower_out(33,50),
			lock_lower_row_in  => s_locks_lower_in(33,50),
			in1                => s_in1(33,50),
			in2                => s_in2(33,50),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(50)
		);
	s_in1(33,50)            <= s_out1(34,50);
	s_in2(33,50)            <= s_out2(34,51);
	s_locks_lower_in(33,50) <= s_locks_lower_out(34,50);

		normal_cell_33_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,51),
			fetch              => s_fetch(33,51),
			data_in            => s_data_in(33,51),
			data_out           => s_data_out(33,51),
			out1               => s_out1(33,51),
			out2               => s_out2(33,51),
			lock_lower_row_out => s_locks_lower_out(33,51),
			lock_lower_row_in  => s_locks_lower_in(33,51),
			in1                => s_in1(33,51),
			in2                => s_in2(33,51),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(51)
		);
	s_in1(33,51)            <= s_out1(34,51);
	s_in2(33,51)            <= s_out2(34,52);
	s_locks_lower_in(33,51) <= s_locks_lower_out(34,51);

		normal_cell_33_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,52),
			fetch              => s_fetch(33,52),
			data_in            => s_data_in(33,52),
			data_out           => s_data_out(33,52),
			out1               => s_out1(33,52),
			out2               => s_out2(33,52),
			lock_lower_row_out => s_locks_lower_out(33,52),
			lock_lower_row_in  => s_locks_lower_in(33,52),
			in1                => s_in1(33,52),
			in2                => s_in2(33,52),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(52)
		);
	s_in1(33,52)            <= s_out1(34,52);
	s_in2(33,52)            <= s_out2(34,53);
	s_locks_lower_in(33,52) <= s_locks_lower_out(34,52);

		normal_cell_33_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,53),
			fetch              => s_fetch(33,53),
			data_in            => s_data_in(33,53),
			data_out           => s_data_out(33,53),
			out1               => s_out1(33,53),
			out2               => s_out2(33,53),
			lock_lower_row_out => s_locks_lower_out(33,53),
			lock_lower_row_in  => s_locks_lower_in(33,53),
			in1                => s_in1(33,53),
			in2                => s_in2(33,53),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(53)
		);
	s_in1(33,53)            <= s_out1(34,53);
	s_in2(33,53)            <= s_out2(34,54);
	s_locks_lower_in(33,53) <= s_locks_lower_out(34,53);

		normal_cell_33_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,54),
			fetch              => s_fetch(33,54),
			data_in            => s_data_in(33,54),
			data_out           => s_data_out(33,54),
			out1               => s_out1(33,54),
			out2               => s_out2(33,54),
			lock_lower_row_out => s_locks_lower_out(33,54),
			lock_lower_row_in  => s_locks_lower_in(33,54),
			in1                => s_in1(33,54),
			in2                => s_in2(33,54),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(54)
		);
	s_in1(33,54)            <= s_out1(34,54);
	s_in2(33,54)            <= s_out2(34,55);
	s_locks_lower_in(33,54) <= s_locks_lower_out(34,54);

		normal_cell_33_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,55),
			fetch              => s_fetch(33,55),
			data_in            => s_data_in(33,55),
			data_out           => s_data_out(33,55),
			out1               => s_out1(33,55),
			out2               => s_out2(33,55),
			lock_lower_row_out => s_locks_lower_out(33,55),
			lock_lower_row_in  => s_locks_lower_in(33,55),
			in1                => s_in1(33,55),
			in2                => s_in2(33,55),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(55)
		);
	s_in1(33,55)            <= s_out1(34,55);
	s_in2(33,55)            <= s_out2(34,56);
	s_locks_lower_in(33,55) <= s_locks_lower_out(34,55);

		normal_cell_33_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,56),
			fetch              => s_fetch(33,56),
			data_in            => s_data_in(33,56),
			data_out           => s_data_out(33,56),
			out1               => s_out1(33,56),
			out2               => s_out2(33,56),
			lock_lower_row_out => s_locks_lower_out(33,56),
			lock_lower_row_in  => s_locks_lower_in(33,56),
			in1                => s_in1(33,56),
			in2                => s_in2(33,56),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(56)
		);
	s_in1(33,56)            <= s_out1(34,56);
	s_in2(33,56)            <= s_out2(34,57);
	s_locks_lower_in(33,56) <= s_locks_lower_out(34,56);

		normal_cell_33_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,57),
			fetch              => s_fetch(33,57),
			data_in            => s_data_in(33,57),
			data_out           => s_data_out(33,57),
			out1               => s_out1(33,57),
			out2               => s_out2(33,57),
			lock_lower_row_out => s_locks_lower_out(33,57),
			lock_lower_row_in  => s_locks_lower_in(33,57),
			in1                => s_in1(33,57),
			in2                => s_in2(33,57),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(57)
		);
	s_in1(33,57)            <= s_out1(34,57);
	s_in2(33,57)            <= s_out2(34,58);
	s_locks_lower_in(33,57) <= s_locks_lower_out(34,57);

		normal_cell_33_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,58),
			fetch              => s_fetch(33,58),
			data_in            => s_data_in(33,58),
			data_out           => s_data_out(33,58),
			out1               => s_out1(33,58),
			out2               => s_out2(33,58),
			lock_lower_row_out => s_locks_lower_out(33,58),
			lock_lower_row_in  => s_locks_lower_in(33,58),
			in1                => s_in1(33,58),
			in2                => s_in2(33,58),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(58)
		);
	s_in1(33,58)            <= s_out1(34,58);
	s_in2(33,58)            <= s_out2(34,59);
	s_locks_lower_in(33,58) <= s_locks_lower_out(34,58);

		normal_cell_33_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,59),
			fetch              => s_fetch(33,59),
			data_in            => s_data_in(33,59),
			data_out           => s_data_out(33,59),
			out1               => s_out1(33,59),
			out2               => s_out2(33,59),
			lock_lower_row_out => s_locks_lower_out(33,59),
			lock_lower_row_in  => s_locks_lower_in(33,59),
			in1                => s_in1(33,59),
			in2                => s_in2(33,59),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(59)
		);
	s_in1(33,59)            <= s_out1(34,59);
	s_in2(33,59)            <= s_out2(34,60);
	s_locks_lower_in(33,59) <= s_locks_lower_out(34,59);

		last_col_cell_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(33,60),
			fetch              => s_fetch(33,60),
			data_in            => s_data_in(33,60),
			data_out           => s_data_out(33,60),
			out1               => s_out1(33,60),
			out2               => s_out2(33,60),
			lock_lower_row_out => s_locks_lower_out(33,60),
			lock_lower_row_in  => s_locks_lower_in(33,60),
			in1                => s_in1(33,60),
			in2                => (others => '0'),
			lock_row           => s_locks(33),
			piv_found          => s_piv_found,
			row_data           => s_row_data(33),
			col_data           => s_col_data(60)
		);
	s_in1(33,60)            <= s_out1(34,60);
	s_locks_lower_in(33,60) <= s_locks_lower_out(34,60);

		normal_cell_34_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,1),
			fetch              => s_fetch(34,1),
			data_in            => s_data_in(34,1),
			data_out           => s_data_out(34,1),
			out1               => s_out1(34,1),
			out2               => s_out2(34,1),
			lock_lower_row_out => s_locks_lower_out(34,1),
			lock_lower_row_in  => s_locks_lower_in(34,1),
			in1                => s_in1(34,1),
			in2                => s_in2(34,1),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(1)
		);
	s_in1(34,1)            <= s_out1(35,1);
	s_in2(34,1)            <= s_out2(35,2);
	s_locks_lower_in(34,1) <= s_locks_lower_out(35,1);

		normal_cell_34_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,2),
			fetch              => s_fetch(34,2),
			data_in            => s_data_in(34,2),
			data_out           => s_data_out(34,2),
			out1               => s_out1(34,2),
			out2               => s_out2(34,2),
			lock_lower_row_out => s_locks_lower_out(34,2),
			lock_lower_row_in  => s_locks_lower_in(34,2),
			in1                => s_in1(34,2),
			in2                => s_in2(34,2),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(2)
		);
	s_in1(34,2)            <= s_out1(35,2);
	s_in2(34,2)            <= s_out2(35,3);
	s_locks_lower_in(34,2) <= s_locks_lower_out(35,2);

		normal_cell_34_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,3),
			fetch              => s_fetch(34,3),
			data_in            => s_data_in(34,3),
			data_out           => s_data_out(34,3),
			out1               => s_out1(34,3),
			out2               => s_out2(34,3),
			lock_lower_row_out => s_locks_lower_out(34,3),
			lock_lower_row_in  => s_locks_lower_in(34,3),
			in1                => s_in1(34,3),
			in2                => s_in2(34,3),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(3)
		);
	s_in1(34,3)            <= s_out1(35,3);
	s_in2(34,3)            <= s_out2(35,4);
	s_locks_lower_in(34,3) <= s_locks_lower_out(35,3);

		normal_cell_34_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,4),
			fetch              => s_fetch(34,4),
			data_in            => s_data_in(34,4),
			data_out           => s_data_out(34,4),
			out1               => s_out1(34,4),
			out2               => s_out2(34,4),
			lock_lower_row_out => s_locks_lower_out(34,4),
			lock_lower_row_in  => s_locks_lower_in(34,4),
			in1                => s_in1(34,4),
			in2                => s_in2(34,4),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(4)
		);
	s_in1(34,4)            <= s_out1(35,4);
	s_in2(34,4)            <= s_out2(35,5);
	s_locks_lower_in(34,4) <= s_locks_lower_out(35,4);

		normal_cell_34_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,5),
			fetch              => s_fetch(34,5),
			data_in            => s_data_in(34,5),
			data_out           => s_data_out(34,5),
			out1               => s_out1(34,5),
			out2               => s_out2(34,5),
			lock_lower_row_out => s_locks_lower_out(34,5),
			lock_lower_row_in  => s_locks_lower_in(34,5),
			in1                => s_in1(34,5),
			in2                => s_in2(34,5),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(5)
		);
	s_in1(34,5)            <= s_out1(35,5);
	s_in2(34,5)            <= s_out2(35,6);
	s_locks_lower_in(34,5) <= s_locks_lower_out(35,5);

		normal_cell_34_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,6),
			fetch              => s_fetch(34,6),
			data_in            => s_data_in(34,6),
			data_out           => s_data_out(34,6),
			out1               => s_out1(34,6),
			out2               => s_out2(34,6),
			lock_lower_row_out => s_locks_lower_out(34,6),
			lock_lower_row_in  => s_locks_lower_in(34,6),
			in1                => s_in1(34,6),
			in2                => s_in2(34,6),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(6)
		);
	s_in1(34,6)            <= s_out1(35,6);
	s_in2(34,6)            <= s_out2(35,7);
	s_locks_lower_in(34,6) <= s_locks_lower_out(35,6);

		normal_cell_34_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,7),
			fetch              => s_fetch(34,7),
			data_in            => s_data_in(34,7),
			data_out           => s_data_out(34,7),
			out1               => s_out1(34,7),
			out2               => s_out2(34,7),
			lock_lower_row_out => s_locks_lower_out(34,7),
			lock_lower_row_in  => s_locks_lower_in(34,7),
			in1                => s_in1(34,7),
			in2                => s_in2(34,7),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(7)
		);
	s_in1(34,7)            <= s_out1(35,7);
	s_in2(34,7)            <= s_out2(35,8);
	s_locks_lower_in(34,7) <= s_locks_lower_out(35,7);

		normal_cell_34_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,8),
			fetch              => s_fetch(34,8),
			data_in            => s_data_in(34,8),
			data_out           => s_data_out(34,8),
			out1               => s_out1(34,8),
			out2               => s_out2(34,8),
			lock_lower_row_out => s_locks_lower_out(34,8),
			lock_lower_row_in  => s_locks_lower_in(34,8),
			in1                => s_in1(34,8),
			in2                => s_in2(34,8),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(8)
		);
	s_in1(34,8)            <= s_out1(35,8);
	s_in2(34,8)            <= s_out2(35,9);
	s_locks_lower_in(34,8) <= s_locks_lower_out(35,8);

		normal_cell_34_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,9),
			fetch              => s_fetch(34,9),
			data_in            => s_data_in(34,9),
			data_out           => s_data_out(34,9),
			out1               => s_out1(34,9),
			out2               => s_out2(34,9),
			lock_lower_row_out => s_locks_lower_out(34,9),
			lock_lower_row_in  => s_locks_lower_in(34,9),
			in1                => s_in1(34,9),
			in2                => s_in2(34,9),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(9)
		);
	s_in1(34,9)            <= s_out1(35,9);
	s_in2(34,9)            <= s_out2(35,10);
	s_locks_lower_in(34,9) <= s_locks_lower_out(35,9);

		normal_cell_34_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,10),
			fetch              => s_fetch(34,10),
			data_in            => s_data_in(34,10),
			data_out           => s_data_out(34,10),
			out1               => s_out1(34,10),
			out2               => s_out2(34,10),
			lock_lower_row_out => s_locks_lower_out(34,10),
			lock_lower_row_in  => s_locks_lower_in(34,10),
			in1                => s_in1(34,10),
			in2                => s_in2(34,10),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(10)
		);
	s_in1(34,10)            <= s_out1(35,10);
	s_in2(34,10)            <= s_out2(35,11);
	s_locks_lower_in(34,10) <= s_locks_lower_out(35,10);

		normal_cell_34_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,11),
			fetch              => s_fetch(34,11),
			data_in            => s_data_in(34,11),
			data_out           => s_data_out(34,11),
			out1               => s_out1(34,11),
			out2               => s_out2(34,11),
			lock_lower_row_out => s_locks_lower_out(34,11),
			lock_lower_row_in  => s_locks_lower_in(34,11),
			in1                => s_in1(34,11),
			in2                => s_in2(34,11),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(11)
		);
	s_in1(34,11)            <= s_out1(35,11);
	s_in2(34,11)            <= s_out2(35,12);
	s_locks_lower_in(34,11) <= s_locks_lower_out(35,11);

		normal_cell_34_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,12),
			fetch              => s_fetch(34,12),
			data_in            => s_data_in(34,12),
			data_out           => s_data_out(34,12),
			out1               => s_out1(34,12),
			out2               => s_out2(34,12),
			lock_lower_row_out => s_locks_lower_out(34,12),
			lock_lower_row_in  => s_locks_lower_in(34,12),
			in1                => s_in1(34,12),
			in2                => s_in2(34,12),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(12)
		);
	s_in1(34,12)            <= s_out1(35,12);
	s_in2(34,12)            <= s_out2(35,13);
	s_locks_lower_in(34,12) <= s_locks_lower_out(35,12);

		normal_cell_34_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,13),
			fetch              => s_fetch(34,13),
			data_in            => s_data_in(34,13),
			data_out           => s_data_out(34,13),
			out1               => s_out1(34,13),
			out2               => s_out2(34,13),
			lock_lower_row_out => s_locks_lower_out(34,13),
			lock_lower_row_in  => s_locks_lower_in(34,13),
			in1                => s_in1(34,13),
			in2                => s_in2(34,13),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(13)
		);
	s_in1(34,13)            <= s_out1(35,13);
	s_in2(34,13)            <= s_out2(35,14);
	s_locks_lower_in(34,13) <= s_locks_lower_out(35,13);

		normal_cell_34_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,14),
			fetch              => s_fetch(34,14),
			data_in            => s_data_in(34,14),
			data_out           => s_data_out(34,14),
			out1               => s_out1(34,14),
			out2               => s_out2(34,14),
			lock_lower_row_out => s_locks_lower_out(34,14),
			lock_lower_row_in  => s_locks_lower_in(34,14),
			in1                => s_in1(34,14),
			in2                => s_in2(34,14),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(14)
		);
	s_in1(34,14)            <= s_out1(35,14);
	s_in2(34,14)            <= s_out2(35,15);
	s_locks_lower_in(34,14) <= s_locks_lower_out(35,14);

		normal_cell_34_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,15),
			fetch              => s_fetch(34,15),
			data_in            => s_data_in(34,15),
			data_out           => s_data_out(34,15),
			out1               => s_out1(34,15),
			out2               => s_out2(34,15),
			lock_lower_row_out => s_locks_lower_out(34,15),
			lock_lower_row_in  => s_locks_lower_in(34,15),
			in1                => s_in1(34,15),
			in2                => s_in2(34,15),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(15)
		);
	s_in1(34,15)            <= s_out1(35,15);
	s_in2(34,15)            <= s_out2(35,16);
	s_locks_lower_in(34,15) <= s_locks_lower_out(35,15);

		normal_cell_34_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,16),
			fetch              => s_fetch(34,16),
			data_in            => s_data_in(34,16),
			data_out           => s_data_out(34,16),
			out1               => s_out1(34,16),
			out2               => s_out2(34,16),
			lock_lower_row_out => s_locks_lower_out(34,16),
			lock_lower_row_in  => s_locks_lower_in(34,16),
			in1                => s_in1(34,16),
			in2                => s_in2(34,16),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(16)
		);
	s_in1(34,16)            <= s_out1(35,16);
	s_in2(34,16)            <= s_out2(35,17);
	s_locks_lower_in(34,16) <= s_locks_lower_out(35,16);

		normal_cell_34_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,17),
			fetch              => s_fetch(34,17),
			data_in            => s_data_in(34,17),
			data_out           => s_data_out(34,17),
			out1               => s_out1(34,17),
			out2               => s_out2(34,17),
			lock_lower_row_out => s_locks_lower_out(34,17),
			lock_lower_row_in  => s_locks_lower_in(34,17),
			in1                => s_in1(34,17),
			in2                => s_in2(34,17),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(17)
		);
	s_in1(34,17)            <= s_out1(35,17);
	s_in2(34,17)            <= s_out2(35,18);
	s_locks_lower_in(34,17) <= s_locks_lower_out(35,17);

		normal_cell_34_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,18),
			fetch              => s_fetch(34,18),
			data_in            => s_data_in(34,18),
			data_out           => s_data_out(34,18),
			out1               => s_out1(34,18),
			out2               => s_out2(34,18),
			lock_lower_row_out => s_locks_lower_out(34,18),
			lock_lower_row_in  => s_locks_lower_in(34,18),
			in1                => s_in1(34,18),
			in2                => s_in2(34,18),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(18)
		);
	s_in1(34,18)            <= s_out1(35,18);
	s_in2(34,18)            <= s_out2(35,19);
	s_locks_lower_in(34,18) <= s_locks_lower_out(35,18);

		normal_cell_34_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,19),
			fetch              => s_fetch(34,19),
			data_in            => s_data_in(34,19),
			data_out           => s_data_out(34,19),
			out1               => s_out1(34,19),
			out2               => s_out2(34,19),
			lock_lower_row_out => s_locks_lower_out(34,19),
			lock_lower_row_in  => s_locks_lower_in(34,19),
			in1                => s_in1(34,19),
			in2                => s_in2(34,19),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(19)
		);
	s_in1(34,19)            <= s_out1(35,19);
	s_in2(34,19)            <= s_out2(35,20);
	s_locks_lower_in(34,19) <= s_locks_lower_out(35,19);

		normal_cell_34_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,20),
			fetch              => s_fetch(34,20),
			data_in            => s_data_in(34,20),
			data_out           => s_data_out(34,20),
			out1               => s_out1(34,20),
			out2               => s_out2(34,20),
			lock_lower_row_out => s_locks_lower_out(34,20),
			lock_lower_row_in  => s_locks_lower_in(34,20),
			in1                => s_in1(34,20),
			in2                => s_in2(34,20),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(20)
		);
	s_in1(34,20)            <= s_out1(35,20);
	s_in2(34,20)            <= s_out2(35,21);
	s_locks_lower_in(34,20) <= s_locks_lower_out(35,20);

		normal_cell_34_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,21),
			fetch              => s_fetch(34,21),
			data_in            => s_data_in(34,21),
			data_out           => s_data_out(34,21),
			out1               => s_out1(34,21),
			out2               => s_out2(34,21),
			lock_lower_row_out => s_locks_lower_out(34,21),
			lock_lower_row_in  => s_locks_lower_in(34,21),
			in1                => s_in1(34,21),
			in2                => s_in2(34,21),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(21)
		);
	s_in1(34,21)            <= s_out1(35,21);
	s_in2(34,21)            <= s_out2(35,22);
	s_locks_lower_in(34,21) <= s_locks_lower_out(35,21);

		normal_cell_34_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,22),
			fetch              => s_fetch(34,22),
			data_in            => s_data_in(34,22),
			data_out           => s_data_out(34,22),
			out1               => s_out1(34,22),
			out2               => s_out2(34,22),
			lock_lower_row_out => s_locks_lower_out(34,22),
			lock_lower_row_in  => s_locks_lower_in(34,22),
			in1                => s_in1(34,22),
			in2                => s_in2(34,22),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(22)
		);
	s_in1(34,22)            <= s_out1(35,22);
	s_in2(34,22)            <= s_out2(35,23);
	s_locks_lower_in(34,22) <= s_locks_lower_out(35,22);

		normal_cell_34_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,23),
			fetch              => s_fetch(34,23),
			data_in            => s_data_in(34,23),
			data_out           => s_data_out(34,23),
			out1               => s_out1(34,23),
			out2               => s_out2(34,23),
			lock_lower_row_out => s_locks_lower_out(34,23),
			lock_lower_row_in  => s_locks_lower_in(34,23),
			in1                => s_in1(34,23),
			in2                => s_in2(34,23),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(23)
		);
	s_in1(34,23)            <= s_out1(35,23);
	s_in2(34,23)            <= s_out2(35,24);
	s_locks_lower_in(34,23) <= s_locks_lower_out(35,23);

		normal_cell_34_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,24),
			fetch              => s_fetch(34,24),
			data_in            => s_data_in(34,24),
			data_out           => s_data_out(34,24),
			out1               => s_out1(34,24),
			out2               => s_out2(34,24),
			lock_lower_row_out => s_locks_lower_out(34,24),
			lock_lower_row_in  => s_locks_lower_in(34,24),
			in1                => s_in1(34,24),
			in2                => s_in2(34,24),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(24)
		);
	s_in1(34,24)            <= s_out1(35,24);
	s_in2(34,24)            <= s_out2(35,25);
	s_locks_lower_in(34,24) <= s_locks_lower_out(35,24);

		normal_cell_34_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,25),
			fetch              => s_fetch(34,25),
			data_in            => s_data_in(34,25),
			data_out           => s_data_out(34,25),
			out1               => s_out1(34,25),
			out2               => s_out2(34,25),
			lock_lower_row_out => s_locks_lower_out(34,25),
			lock_lower_row_in  => s_locks_lower_in(34,25),
			in1                => s_in1(34,25),
			in2                => s_in2(34,25),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(25)
		);
	s_in1(34,25)            <= s_out1(35,25);
	s_in2(34,25)            <= s_out2(35,26);
	s_locks_lower_in(34,25) <= s_locks_lower_out(35,25);

		normal_cell_34_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,26),
			fetch              => s_fetch(34,26),
			data_in            => s_data_in(34,26),
			data_out           => s_data_out(34,26),
			out1               => s_out1(34,26),
			out2               => s_out2(34,26),
			lock_lower_row_out => s_locks_lower_out(34,26),
			lock_lower_row_in  => s_locks_lower_in(34,26),
			in1                => s_in1(34,26),
			in2                => s_in2(34,26),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(26)
		);
	s_in1(34,26)            <= s_out1(35,26);
	s_in2(34,26)            <= s_out2(35,27);
	s_locks_lower_in(34,26) <= s_locks_lower_out(35,26);

		normal_cell_34_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,27),
			fetch              => s_fetch(34,27),
			data_in            => s_data_in(34,27),
			data_out           => s_data_out(34,27),
			out1               => s_out1(34,27),
			out2               => s_out2(34,27),
			lock_lower_row_out => s_locks_lower_out(34,27),
			lock_lower_row_in  => s_locks_lower_in(34,27),
			in1                => s_in1(34,27),
			in2                => s_in2(34,27),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(27)
		);
	s_in1(34,27)            <= s_out1(35,27);
	s_in2(34,27)            <= s_out2(35,28);
	s_locks_lower_in(34,27) <= s_locks_lower_out(35,27);

		normal_cell_34_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,28),
			fetch              => s_fetch(34,28),
			data_in            => s_data_in(34,28),
			data_out           => s_data_out(34,28),
			out1               => s_out1(34,28),
			out2               => s_out2(34,28),
			lock_lower_row_out => s_locks_lower_out(34,28),
			lock_lower_row_in  => s_locks_lower_in(34,28),
			in1                => s_in1(34,28),
			in2                => s_in2(34,28),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(28)
		);
	s_in1(34,28)            <= s_out1(35,28);
	s_in2(34,28)            <= s_out2(35,29);
	s_locks_lower_in(34,28) <= s_locks_lower_out(35,28);

		normal_cell_34_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,29),
			fetch              => s_fetch(34,29),
			data_in            => s_data_in(34,29),
			data_out           => s_data_out(34,29),
			out1               => s_out1(34,29),
			out2               => s_out2(34,29),
			lock_lower_row_out => s_locks_lower_out(34,29),
			lock_lower_row_in  => s_locks_lower_in(34,29),
			in1                => s_in1(34,29),
			in2                => s_in2(34,29),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(29)
		);
	s_in1(34,29)            <= s_out1(35,29);
	s_in2(34,29)            <= s_out2(35,30);
	s_locks_lower_in(34,29) <= s_locks_lower_out(35,29);

		normal_cell_34_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,30),
			fetch              => s_fetch(34,30),
			data_in            => s_data_in(34,30),
			data_out           => s_data_out(34,30),
			out1               => s_out1(34,30),
			out2               => s_out2(34,30),
			lock_lower_row_out => s_locks_lower_out(34,30),
			lock_lower_row_in  => s_locks_lower_in(34,30),
			in1                => s_in1(34,30),
			in2                => s_in2(34,30),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(30)
		);
	s_in1(34,30)            <= s_out1(35,30);
	s_in2(34,30)            <= s_out2(35,31);
	s_locks_lower_in(34,30) <= s_locks_lower_out(35,30);

		normal_cell_34_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,31),
			fetch              => s_fetch(34,31),
			data_in            => s_data_in(34,31),
			data_out           => s_data_out(34,31),
			out1               => s_out1(34,31),
			out2               => s_out2(34,31),
			lock_lower_row_out => s_locks_lower_out(34,31),
			lock_lower_row_in  => s_locks_lower_in(34,31),
			in1                => s_in1(34,31),
			in2                => s_in2(34,31),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(31)
		);
	s_in1(34,31)            <= s_out1(35,31);
	s_in2(34,31)            <= s_out2(35,32);
	s_locks_lower_in(34,31) <= s_locks_lower_out(35,31);

		normal_cell_34_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,32),
			fetch              => s_fetch(34,32),
			data_in            => s_data_in(34,32),
			data_out           => s_data_out(34,32),
			out1               => s_out1(34,32),
			out2               => s_out2(34,32),
			lock_lower_row_out => s_locks_lower_out(34,32),
			lock_lower_row_in  => s_locks_lower_in(34,32),
			in1                => s_in1(34,32),
			in2                => s_in2(34,32),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(32)
		);
	s_in1(34,32)            <= s_out1(35,32);
	s_in2(34,32)            <= s_out2(35,33);
	s_locks_lower_in(34,32) <= s_locks_lower_out(35,32);

		normal_cell_34_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,33),
			fetch              => s_fetch(34,33),
			data_in            => s_data_in(34,33),
			data_out           => s_data_out(34,33),
			out1               => s_out1(34,33),
			out2               => s_out2(34,33),
			lock_lower_row_out => s_locks_lower_out(34,33),
			lock_lower_row_in  => s_locks_lower_in(34,33),
			in1                => s_in1(34,33),
			in2                => s_in2(34,33),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(33)
		);
	s_in1(34,33)            <= s_out1(35,33);
	s_in2(34,33)            <= s_out2(35,34);
	s_locks_lower_in(34,33) <= s_locks_lower_out(35,33);

		normal_cell_34_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,34),
			fetch              => s_fetch(34,34),
			data_in            => s_data_in(34,34),
			data_out           => s_data_out(34,34),
			out1               => s_out1(34,34),
			out2               => s_out2(34,34),
			lock_lower_row_out => s_locks_lower_out(34,34),
			lock_lower_row_in  => s_locks_lower_in(34,34),
			in1                => s_in1(34,34),
			in2                => s_in2(34,34),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(34)
		);
	s_in1(34,34)            <= s_out1(35,34);
	s_in2(34,34)            <= s_out2(35,35);
	s_locks_lower_in(34,34) <= s_locks_lower_out(35,34);

		normal_cell_34_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,35),
			fetch              => s_fetch(34,35),
			data_in            => s_data_in(34,35),
			data_out           => s_data_out(34,35),
			out1               => s_out1(34,35),
			out2               => s_out2(34,35),
			lock_lower_row_out => s_locks_lower_out(34,35),
			lock_lower_row_in  => s_locks_lower_in(34,35),
			in1                => s_in1(34,35),
			in2                => s_in2(34,35),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(35)
		);
	s_in1(34,35)            <= s_out1(35,35);
	s_in2(34,35)            <= s_out2(35,36);
	s_locks_lower_in(34,35) <= s_locks_lower_out(35,35);

		normal_cell_34_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,36),
			fetch              => s_fetch(34,36),
			data_in            => s_data_in(34,36),
			data_out           => s_data_out(34,36),
			out1               => s_out1(34,36),
			out2               => s_out2(34,36),
			lock_lower_row_out => s_locks_lower_out(34,36),
			lock_lower_row_in  => s_locks_lower_in(34,36),
			in1                => s_in1(34,36),
			in2                => s_in2(34,36),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(36)
		);
	s_in1(34,36)            <= s_out1(35,36);
	s_in2(34,36)            <= s_out2(35,37);
	s_locks_lower_in(34,36) <= s_locks_lower_out(35,36);

		normal_cell_34_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,37),
			fetch              => s_fetch(34,37),
			data_in            => s_data_in(34,37),
			data_out           => s_data_out(34,37),
			out1               => s_out1(34,37),
			out2               => s_out2(34,37),
			lock_lower_row_out => s_locks_lower_out(34,37),
			lock_lower_row_in  => s_locks_lower_in(34,37),
			in1                => s_in1(34,37),
			in2                => s_in2(34,37),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(37)
		);
	s_in1(34,37)            <= s_out1(35,37);
	s_in2(34,37)            <= s_out2(35,38);
	s_locks_lower_in(34,37) <= s_locks_lower_out(35,37);

		normal_cell_34_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,38),
			fetch              => s_fetch(34,38),
			data_in            => s_data_in(34,38),
			data_out           => s_data_out(34,38),
			out1               => s_out1(34,38),
			out2               => s_out2(34,38),
			lock_lower_row_out => s_locks_lower_out(34,38),
			lock_lower_row_in  => s_locks_lower_in(34,38),
			in1                => s_in1(34,38),
			in2                => s_in2(34,38),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(38)
		);
	s_in1(34,38)            <= s_out1(35,38);
	s_in2(34,38)            <= s_out2(35,39);
	s_locks_lower_in(34,38) <= s_locks_lower_out(35,38);

		normal_cell_34_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,39),
			fetch              => s_fetch(34,39),
			data_in            => s_data_in(34,39),
			data_out           => s_data_out(34,39),
			out1               => s_out1(34,39),
			out2               => s_out2(34,39),
			lock_lower_row_out => s_locks_lower_out(34,39),
			lock_lower_row_in  => s_locks_lower_in(34,39),
			in1                => s_in1(34,39),
			in2                => s_in2(34,39),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(39)
		);
	s_in1(34,39)            <= s_out1(35,39);
	s_in2(34,39)            <= s_out2(35,40);
	s_locks_lower_in(34,39) <= s_locks_lower_out(35,39);

		normal_cell_34_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,40),
			fetch              => s_fetch(34,40),
			data_in            => s_data_in(34,40),
			data_out           => s_data_out(34,40),
			out1               => s_out1(34,40),
			out2               => s_out2(34,40),
			lock_lower_row_out => s_locks_lower_out(34,40),
			lock_lower_row_in  => s_locks_lower_in(34,40),
			in1                => s_in1(34,40),
			in2                => s_in2(34,40),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(40)
		);
	s_in1(34,40)            <= s_out1(35,40);
	s_in2(34,40)            <= s_out2(35,41);
	s_locks_lower_in(34,40) <= s_locks_lower_out(35,40);

		normal_cell_34_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,41),
			fetch              => s_fetch(34,41),
			data_in            => s_data_in(34,41),
			data_out           => s_data_out(34,41),
			out1               => s_out1(34,41),
			out2               => s_out2(34,41),
			lock_lower_row_out => s_locks_lower_out(34,41),
			lock_lower_row_in  => s_locks_lower_in(34,41),
			in1                => s_in1(34,41),
			in2                => s_in2(34,41),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(41)
		);
	s_in1(34,41)            <= s_out1(35,41);
	s_in2(34,41)            <= s_out2(35,42);
	s_locks_lower_in(34,41) <= s_locks_lower_out(35,41);

		normal_cell_34_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,42),
			fetch              => s_fetch(34,42),
			data_in            => s_data_in(34,42),
			data_out           => s_data_out(34,42),
			out1               => s_out1(34,42),
			out2               => s_out2(34,42),
			lock_lower_row_out => s_locks_lower_out(34,42),
			lock_lower_row_in  => s_locks_lower_in(34,42),
			in1                => s_in1(34,42),
			in2                => s_in2(34,42),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(42)
		);
	s_in1(34,42)            <= s_out1(35,42);
	s_in2(34,42)            <= s_out2(35,43);
	s_locks_lower_in(34,42) <= s_locks_lower_out(35,42);

		normal_cell_34_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,43),
			fetch              => s_fetch(34,43),
			data_in            => s_data_in(34,43),
			data_out           => s_data_out(34,43),
			out1               => s_out1(34,43),
			out2               => s_out2(34,43),
			lock_lower_row_out => s_locks_lower_out(34,43),
			lock_lower_row_in  => s_locks_lower_in(34,43),
			in1                => s_in1(34,43),
			in2                => s_in2(34,43),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(43)
		);
	s_in1(34,43)            <= s_out1(35,43);
	s_in2(34,43)            <= s_out2(35,44);
	s_locks_lower_in(34,43) <= s_locks_lower_out(35,43);

		normal_cell_34_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,44),
			fetch              => s_fetch(34,44),
			data_in            => s_data_in(34,44),
			data_out           => s_data_out(34,44),
			out1               => s_out1(34,44),
			out2               => s_out2(34,44),
			lock_lower_row_out => s_locks_lower_out(34,44),
			lock_lower_row_in  => s_locks_lower_in(34,44),
			in1                => s_in1(34,44),
			in2                => s_in2(34,44),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(44)
		);
	s_in1(34,44)            <= s_out1(35,44);
	s_in2(34,44)            <= s_out2(35,45);
	s_locks_lower_in(34,44) <= s_locks_lower_out(35,44);

		normal_cell_34_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,45),
			fetch              => s_fetch(34,45),
			data_in            => s_data_in(34,45),
			data_out           => s_data_out(34,45),
			out1               => s_out1(34,45),
			out2               => s_out2(34,45),
			lock_lower_row_out => s_locks_lower_out(34,45),
			lock_lower_row_in  => s_locks_lower_in(34,45),
			in1                => s_in1(34,45),
			in2                => s_in2(34,45),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(45)
		);
	s_in1(34,45)            <= s_out1(35,45);
	s_in2(34,45)            <= s_out2(35,46);
	s_locks_lower_in(34,45) <= s_locks_lower_out(35,45);

		normal_cell_34_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,46),
			fetch              => s_fetch(34,46),
			data_in            => s_data_in(34,46),
			data_out           => s_data_out(34,46),
			out1               => s_out1(34,46),
			out2               => s_out2(34,46),
			lock_lower_row_out => s_locks_lower_out(34,46),
			lock_lower_row_in  => s_locks_lower_in(34,46),
			in1                => s_in1(34,46),
			in2                => s_in2(34,46),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(46)
		);
	s_in1(34,46)            <= s_out1(35,46);
	s_in2(34,46)            <= s_out2(35,47);
	s_locks_lower_in(34,46) <= s_locks_lower_out(35,46);

		normal_cell_34_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,47),
			fetch              => s_fetch(34,47),
			data_in            => s_data_in(34,47),
			data_out           => s_data_out(34,47),
			out1               => s_out1(34,47),
			out2               => s_out2(34,47),
			lock_lower_row_out => s_locks_lower_out(34,47),
			lock_lower_row_in  => s_locks_lower_in(34,47),
			in1                => s_in1(34,47),
			in2                => s_in2(34,47),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(47)
		);
	s_in1(34,47)            <= s_out1(35,47);
	s_in2(34,47)            <= s_out2(35,48);
	s_locks_lower_in(34,47) <= s_locks_lower_out(35,47);

		normal_cell_34_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,48),
			fetch              => s_fetch(34,48),
			data_in            => s_data_in(34,48),
			data_out           => s_data_out(34,48),
			out1               => s_out1(34,48),
			out2               => s_out2(34,48),
			lock_lower_row_out => s_locks_lower_out(34,48),
			lock_lower_row_in  => s_locks_lower_in(34,48),
			in1                => s_in1(34,48),
			in2                => s_in2(34,48),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(48)
		);
	s_in1(34,48)            <= s_out1(35,48);
	s_in2(34,48)            <= s_out2(35,49);
	s_locks_lower_in(34,48) <= s_locks_lower_out(35,48);

		normal_cell_34_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,49),
			fetch              => s_fetch(34,49),
			data_in            => s_data_in(34,49),
			data_out           => s_data_out(34,49),
			out1               => s_out1(34,49),
			out2               => s_out2(34,49),
			lock_lower_row_out => s_locks_lower_out(34,49),
			lock_lower_row_in  => s_locks_lower_in(34,49),
			in1                => s_in1(34,49),
			in2                => s_in2(34,49),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(49)
		);
	s_in1(34,49)            <= s_out1(35,49);
	s_in2(34,49)            <= s_out2(35,50);
	s_locks_lower_in(34,49) <= s_locks_lower_out(35,49);

		normal_cell_34_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,50),
			fetch              => s_fetch(34,50),
			data_in            => s_data_in(34,50),
			data_out           => s_data_out(34,50),
			out1               => s_out1(34,50),
			out2               => s_out2(34,50),
			lock_lower_row_out => s_locks_lower_out(34,50),
			lock_lower_row_in  => s_locks_lower_in(34,50),
			in1                => s_in1(34,50),
			in2                => s_in2(34,50),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(50)
		);
	s_in1(34,50)            <= s_out1(35,50);
	s_in2(34,50)            <= s_out2(35,51);
	s_locks_lower_in(34,50) <= s_locks_lower_out(35,50);

		normal_cell_34_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,51),
			fetch              => s_fetch(34,51),
			data_in            => s_data_in(34,51),
			data_out           => s_data_out(34,51),
			out1               => s_out1(34,51),
			out2               => s_out2(34,51),
			lock_lower_row_out => s_locks_lower_out(34,51),
			lock_lower_row_in  => s_locks_lower_in(34,51),
			in1                => s_in1(34,51),
			in2                => s_in2(34,51),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(51)
		);
	s_in1(34,51)            <= s_out1(35,51);
	s_in2(34,51)            <= s_out2(35,52);
	s_locks_lower_in(34,51) <= s_locks_lower_out(35,51);

		normal_cell_34_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,52),
			fetch              => s_fetch(34,52),
			data_in            => s_data_in(34,52),
			data_out           => s_data_out(34,52),
			out1               => s_out1(34,52),
			out2               => s_out2(34,52),
			lock_lower_row_out => s_locks_lower_out(34,52),
			lock_lower_row_in  => s_locks_lower_in(34,52),
			in1                => s_in1(34,52),
			in2                => s_in2(34,52),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(52)
		);
	s_in1(34,52)            <= s_out1(35,52);
	s_in2(34,52)            <= s_out2(35,53);
	s_locks_lower_in(34,52) <= s_locks_lower_out(35,52);

		normal_cell_34_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,53),
			fetch              => s_fetch(34,53),
			data_in            => s_data_in(34,53),
			data_out           => s_data_out(34,53),
			out1               => s_out1(34,53),
			out2               => s_out2(34,53),
			lock_lower_row_out => s_locks_lower_out(34,53),
			lock_lower_row_in  => s_locks_lower_in(34,53),
			in1                => s_in1(34,53),
			in2                => s_in2(34,53),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(53)
		);
	s_in1(34,53)            <= s_out1(35,53);
	s_in2(34,53)            <= s_out2(35,54);
	s_locks_lower_in(34,53) <= s_locks_lower_out(35,53);

		normal_cell_34_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,54),
			fetch              => s_fetch(34,54),
			data_in            => s_data_in(34,54),
			data_out           => s_data_out(34,54),
			out1               => s_out1(34,54),
			out2               => s_out2(34,54),
			lock_lower_row_out => s_locks_lower_out(34,54),
			lock_lower_row_in  => s_locks_lower_in(34,54),
			in1                => s_in1(34,54),
			in2                => s_in2(34,54),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(54)
		);
	s_in1(34,54)            <= s_out1(35,54);
	s_in2(34,54)            <= s_out2(35,55);
	s_locks_lower_in(34,54) <= s_locks_lower_out(35,54);

		normal_cell_34_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,55),
			fetch              => s_fetch(34,55),
			data_in            => s_data_in(34,55),
			data_out           => s_data_out(34,55),
			out1               => s_out1(34,55),
			out2               => s_out2(34,55),
			lock_lower_row_out => s_locks_lower_out(34,55),
			lock_lower_row_in  => s_locks_lower_in(34,55),
			in1                => s_in1(34,55),
			in2                => s_in2(34,55),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(55)
		);
	s_in1(34,55)            <= s_out1(35,55);
	s_in2(34,55)            <= s_out2(35,56);
	s_locks_lower_in(34,55) <= s_locks_lower_out(35,55);

		normal_cell_34_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,56),
			fetch              => s_fetch(34,56),
			data_in            => s_data_in(34,56),
			data_out           => s_data_out(34,56),
			out1               => s_out1(34,56),
			out2               => s_out2(34,56),
			lock_lower_row_out => s_locks_lower_out(34,56),
			lock_lower_row_in  => s_locks_lower_in(34,56),
			in1                => s_in1(34,56),
			in2                => s_in2(34,56),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(56)
		);
	s_in1(34,56)            <= s_out1(35,56);
	s_in2(34,56)            <= s_out2(35,57);
	s_locks_lower_in(34,56) <= s_locks_lower_out(35,56);

		normal_cell_34_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,57),
			fetch              => s_fetch(34,57),
			data_in            => s_data_in(34,57),
			data_out           => s_data_out(34,57),
			out1               => s_out1(34,57),
			out2               => s_out2(34,57),
			lock_lower_row_out => s_locks_lower_out(34,57),
			lock_lower_row_in  => s_locks_lower_in(34,57),
			in1                => s_in1(34,57),
			in2                => s_in2(34,57),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(57)
		);
	s_in1(34,57)            <= s_out1(35,57);
	s_in2(34,57)            <= s_out2(35,58);
	s_locks_lower_in(34,57) <= s_locks_lower_out(35,57);

		normal_cell_34_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,58),
			fetch              => s_fetch(34,58),
			data_in            => s_data_in(34,58),
			data_out           => s_data_out(34,58),
			out1               => s_out1(34,58),
			out2               => s_out2(34,58),
			lock_lower_row_out => s_locks_lower_out(34,58),
			lock_lower_row_in  => s_locks_lower_in(34,58),
			in1                => s_in1(34,58),
			in2                => s_in2(34,58),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(58)
		);
	s_in1(34,58)            <= s_out1(35,58);
	s_in2(34,58)            <= s_out2(35,59);
	s_locks_lower_in(34,58) <= s_locks_lower_out(35,58);

		normal_cell_34_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,59),
			fetch              => s_fetch(34,59),
			data_in            => s_data_in(34,59),
			data_out           => s_data_out(34,59),
			out1               => s_out1(34,59),
			out2               => s_out2(34,59),
			lock_lower_row_out => s_locks_lower_out(34,59),
			lock_lower_row_in  => s_locks_lower_in(34,59),
			in1                => s_in1(34,59),
			in2                => s_in2(34,59),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(59)
		);
	s_in1(34,59)            <= s_out1(35,59);
	s_in2(34,59)            <= s_out2(35,60);
	s_locks_lower_in(34,59) <= s_locks_lower_out(35,59);

		last_col_cell_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(34,60),
			fetch              => s_fetch(34,60),
			data_in            => s_data_in(34,60),
			data_out           => s_data_out(34,60),
			out1               => s_out1(34,60),
			out2               => s_out2(34,60),
			lock_lower_row_out => s_locks_lower_out(34,60),
			lock_lower_row_in  => s_locks_lower_in(34,60),
			in1                => s_in1(34,60),
			in2                => (others => '0'),
			lock_row           => s_locks(34),
			piv_found          => s_piv_found,
			row_data           => s_row_data(34),
			col_data           => s_col_data(60)
		);
	s_in1(34,60)            <= s_out1(35,60);
	s_locks_lower_in(34,60) <= s_locks_lower_out(35,60);

		normal_cell_35_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,1),
			fetch              => s_fetch(35,1),
			data_in            => s_data_in(35,1),
			data_out           => s_data_out(35,1),
			out1               => s_out1(35,1),
			out2               => s_out2(35,1),
			lock_lower_row_out => s_locks_lower_out(35,1),
			lock_lower_row_in  => s_locks_lower_in(35,1),
			in1                => s_in1(35,1),
			in2                => s_in2(35,1),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(1)
		);
	s_in1(35,1)            <= s_out1(36,1);
	s_in2(35,1)            <= s_out2(36,2);
	s_locks_lower_in(35,1) <= s_locks_lower_out(36,1);

		normal_cell_35_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,2),
			fetch              => s_fetch(35,2),
			data_in            => s_data_in(35,2),
			data_out           => s_data_out(35,2),
			out1               => s_out1(35,2),
			out2               => s_out2(35,2),
			lock_lower_row_out => s_locks_lower_out(35,2),
			lock_lower_row_in  => s_locks_lower_in(35,2),
			in1                => s_in1(35,2),
			in2                => s_in2(35,2),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(2)
		);
	s_in1(35,2)            <= s_out1(36,2);
	s_in2(35,2)            <= s_out2(36,3);
	s_locks_lower_in(35,2) <= s_locks_lower_out(36,2);

		normal_cell_35_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,3),
			fetch              => s_fetch(35,3),
			data_in            => s_data_in(35,3),
			data_out           => s_data_out(35,3),
			out1               => s_out1(35,3),
			out2               => s_out2(35,3),
			lock_lower_row_out => s_locks_lower_out(35,3),
			lock_lower_row_in  => s_locks_lower_in(35,3),
			in1                => s_in1(35,3),
			in2                => s_in2(35,3),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(3)
		);
	s_in1(35,3)            <= s_out1(36,3);
	s_in2(35,3)            <= s_out2(36,4);
	s_locks_lower_in(35,3) <= s_locks_lower_out(36,3);

		normal_cell_35_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,4),
			fetch              => s_fetch(35,4),
			data_in            => s_data_in(35,4),
			data_out           => s_data_out(35,4),
			out1               => s_out1(35,4),
			out2               => s_out2(35,4),
			lock_lower_row_out => s_locks_lower_out(35,4),
			lock_lower_row_in  => s_locks_lower_in(35,4),
			in1                => s_in1(35,4),
			in2                => s_in2(35,4),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(4)
		);
	s_in1(35,4)            <= s_out1(36,4);
	s_in2(35,4)            <= s_out2(36,5);
	s_locks_lower_in(35,4) <= s_locks_lower_out(36,4);

		normal_cell_35_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,5),
			fetch              => s_fetch(35,5),
			data_in            => s_data_in(35,5),
			data_out           => s_data_out(35,5),
			out1               => s_out1(35,5),
			out2               => s_out2(35,5),
			lock_lower_row_out => s_locks_lower_out(35,5),
			lock_lower_row_in  => s_locks_lower_in(35,5),
			in1                => s_in1(35,5),
			in2                => s_in2(35,5),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(5)
		);
	s_in1(35,5)            <= s_out1(36,5);
	s_in2(35,5)            <= s_out2(36,6);
	s_locks_lower_in(35,5) <= s_locks_lower_out(36,5);

		normal_cell_35_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,6),
			fetch              => s_fetch(35,6),
			data_in            => s_data_in(35,6),
			data_out           => s_data_out(35,6),
			out1               => s_out1(35,6),
			out2               => s_out2(35,6),
			lock_lower_row_out => s_locks_lower_out(35,6),
			lock_lower_row_in  => s_locks_lower_in(35,6),
			in1                => s_in1(35,6),
			in2                => s_in2(35,6),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(6)
		);
	s_in1(35,6)            <= s_out1(36,6);
	s_in2(35,6)            <= s_out2(36,7);
	s_locks_lower_in(35,6) <= s_locks_lower_out(36,6);

		normal_cell_35_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,7),
			fetch              => s_fetch(35,7),
			data_in            => s_data_in(35,7),
			data_out           => s_data_out(35,7),
			out1               => s_out1(35,7),
			out2               => s_out2(35,7),
			lock_lower_row_out => s_locks_lower_out(35,7),
			lock_lower_row_in  => s_locks_lower_in(35,7),
			in1                => s_in1(35,7),
			in2                => s_in2(35,7),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(7)
		);
	s_in1(35,7)            <= s_out1(36,7);
	s_in2(35,7)            <= s_out2(36,8);
	s_locks_lower_in(35,7) <= s_locks_lower_out(36,7);

		normal_cell_35_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,8),
			fetch              => s_fetch(35,8),
			data_in            => s_data_in(35,8),
			data_out           => s_data_out(35,8),
			out1               => s_out1(35,8),
			out2               => s_out2(35,8),
			lock_lower_row_out => s_locks_lower_out(35,8),
			lock_lower_row_in  => s_locks_lower_in(35,8),
			in1                => s_in1(35,8),
			in2                => s_in2(35,8),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(8)
		);
	s_in1(35,8)            <= s_out1(36,8);
	s_in2(35,8)            <= s_out2(36,9);
	s_locks_lower_in(35,8) <= s_locks_lower_out(36,8);

		normal_cell_35_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,9),
			fetch              => s_fetch(35,9),
			data_in            => s_data_in(35,9),
			data_out           => s_data_out(35,9),
			out1               => s_out1(35,9),
			out2               => s_out2(35,9),
			lock_lower_row_out => s_locks_lower_out(35,9),
			lock_lower_row_in  => s_locks_lower_in(35,9),
			in1                => s_in1(35,9),
			in2                => s_in2(35,9),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(9)
		);
	s_in1(35,9)            <= s_out1(36,9);
	s_in2(35,9)            <= s_out2(36,10);
	s_locks_lower_in(35,9) <= s_locks_lower_out(36,9);

		normal_cell_35_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,10),
			fetch              => s_fetch(35,10),
			data_in            => s_data_in(35,10),
			data_out           => s_data_out(35,10),
			out1               => s_out1(35,10),
			out2               => s_out2(35,10),
			lock_lower_row_out => s_locks_lower_out(35,10),
			lock_lower_row_in  => s_locks_lower_in(35,10),
			in1                => s_in1(35,10),
			in2                => s_in2(35,10),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(10)
		);
	s_in1(35,10)            <= s_out1(36,10);
	s_in2(35,10)            <= s_out2(36,11);
	s_locks_lower_in(35,10) <= s_locks_lower_out(36,10);

		normal_cell_35_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,11),
			fetch              => s_fetch(35,11),
			data_in            => s_data_in(35,11),
			data_out           => s_data_out(35,11),
			out1               => s_out1(35,11),
			out2               => s_out2(35,11),
			lock_lower_row_out => s_locks_lower_out(35,11),
			lock_lower_row_in  => s_locks_lower_in(35,11),
			in1                => s_in1(35,11),
			in2                => s_in2(35,11),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(11)
		);
	s_in1(35,11)            <= s_out1(36,11);
	s_in2(35,11)            <= s_out2(36,12);
	s_locks_lower_in(35,11) <= s_locks_lower_out(36,11);

		normal_cell_35_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,12),
			fetch              => s_fetch(35,12),
			data_in            => s_data_in(35,12),
			data_out           => s_data_out(35,12),
			out1               => s_out1(35,12),
			out2               => s_out2(35,12),
			lock_lower_row_out => s_locks_lower_out(35,12),
			lock_lower_row_in  => s_locks_lower_in(35,12),
			in1                => s_in1(35,12),
			in2                => s_in2(35,12),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(12)
		);
	s_in1(35,12)            <= s_out1(36,12);
	s_in2(35,12)            <= s_out2(36,13);
	s_locks_lower_in(35,12) <= s_locks_lower_out(36,12);

		normal_cell_35_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,13),
			fetch              => s_fetch(35,13),
			data_in            => s_data_in(35,13),
			data_out           => s_data_out(35,13),
			out1               => s_out1(35,13),
			out2               => s_out2(35,13),
			lock_lower_row_out => s_locks_lower_out(35,13),
			lock_lower_row_in  => s_locks_lower_in(35,13),
			in1                => s_in1(35,13),
			in2                => s_in2(35,13),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(13)
		);
	s_in1(35,13)            <= s_out1(36,13);
	s_in2(35,13)            <= s_out2(36,14);
	s_locks_lower_in(35,13) <= s_locks_lower_out(36,13);

		normal_cell_35_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,14),
			fetch              => s_fetch(35,14),
			data_in            => s_data_in(35,14),
			data_out           => s_data_out(35,14),
			out1               => s_out1(35,14),
			out2               => s_out2(35,14),
			lock_lower_row_out => s_locks_lower_out(35,14),
			lock_lower_row_in  => s_locks_lower_in(35,14),
			in1                => s_in1(35,14),
			in2                => s_in2(35,14),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(14)
		);
	s_in1(35,14)            <= s_out1(36,14);
	s_in2(35,14)            <= s_out2(36,15);
	s_locks_lower_in(35,14) <= s_locks_lower_out(36,14);

		normal_cell_35_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,15),
			fetch              => s_fetch(35,15),
			data_in            => s_data_in(35,15),
			data_out           => s_data_out(35,15),
			out1               => s_out1(35,15),
			out2               => s_out2(35,15),
			lock_lower_row_out => s_locks_lower_out(35,15),
			lock_lower_row_in  => s_locks_lower_in(35,15),
			in1                => s_in1(35,15),
			in2                => s_in2(35,15),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(15)
		);
	s_in1(35,15)            <= s_out1(36,15);
	s_in2(35,15)            <= s_out2(36,16);
	s_locks_lower_in(35,15) <= s_locks_lower_out(36,15);

		normal_cell_35_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,16),
			fetch              => s_fetch(35,16),
			data_in            => s_data_in(35,16),
			data_out           => s_data_out(35,16),
			out1               => s_out1(35,16),
			out2               => s_out2(35,16),
			lock_lower_row_out => s_locks_lower_out(35,16),
			lock_lower_row_in  => s_locks_lower_in(35,16),
			in1                => s_in1(35,16),
			in2                => s_in2(35,16),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(16)
		);
	s_in1(35,16)            <= s_out1(36,16);
	s_in2(35,16)            <= s_out2(36,17);
	s_locks_lower_in(35,16) <= s_locks_lower_out(36,16);

		normal_cell_35_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,17),
			fetch              => s_fetch(35,17),
			data_in            => s_data_in(35,17),
			data_out           => s_data_out(35,17),
			out1               => s_out1(35,17),
			out2               => s_out2(35,17),
			lock_lower_row_out => s_locks_lower_out(35,17),
			lock_lower_row_in  => s_locks_lower_in(35,17),
			in1                => s_in1(35,17),
			in2                => s_in2(35,17),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(17)
		);
	s_in1(35,17)            <= s_out1(36,17);
	s_in2(35,17)            <= s_out2(36,18);
	s_locks_lower_in(35,17) <= s_locks_lower_out(36,17);

		normal_cell_35_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,18),
			fetch              => s_fetch(35,18),
			data_in            => s_data_in(35,18),
			data_out           => s_data_out(35,18),
			out1               => s_out1(35,18),
			out2               => s_out2(35,18),
			lock_lower_row_out => s_locks_lower_out(35,18),
			lock_lower_row_in  => s_locks_lower_in(35,18),
			in1                => s_in1(35,18),
			in2                => s_in2(35,18),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(18)
		);
	s_in1(35,18)            <= s_out1(36,18);
	s_in2(35,18)            <= s_out2(36,19);
	s_locks_lower_in(35,18) <= s_locks_lower_out(36,18);

		normal_cell_35_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,19),
			fetch              => s_fetch(35,19),
			data_in            => s_data_in(35,19),
			data_out           => s_data_out(35,19),
			out1               => s_out1(35,19),
			out2               => s_out2(35,19),
			lock_lower_row_out => s_locks_lower_out(35,19),
			lock_lower_row_in  => s_locks_lower_in(35,19),
			in1                => s_in1(35,19),
			in2                => s_in2(35,19),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(19)
		);
	s_in1(35,19)            <= s_out1(36,19);
	s_in2(35,19)            <= s_out2(36,20);
	s_locks_lower_in(35,19) <= s_locks_lower_out(36,19);

		normal_cell_35_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,20),
			fetch              => s_fetch(35,20),
			data_in            => s_data_in(35,20),
			data_out           => s_data_out(35,20),
			out1               => s_out1(35,20),
			out2               => s_out2(35,20),
			lock_lower_row_out => s_locks_lower_out(35,20),
			lock_lower_row_in  => s_locks_lower_in(35,20),
			in1                => s_in1(35,20),
			in2                => s_in2(35,20),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(20)
		);
	s_in1(35,20)            <= s_out1(36,20);
	s_in2(35,20)            <= s_out2(36,21);
	s_locks_lower_in(35,20) <= s_locks_lower_out(36,20);

		normal_cell_35_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,21),
			fetch              => s_fetch(35,21),
			data_in            => s_data_in(35,21),
			data_out           => s_data_out(35,21),
			out1               => s_out1(35,21),
			out2               => s_out2(35,21),
			lock_lower_row_out => s_locks_lower_out(35,21),
			lock_lower_row_in  => s_locks_lower_in(35,21),
			in1                => s_in1(35,21),
			in2                => s_in2(35,21),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(21)
		);
	s_in1(35,21)            <= s_out1(36,21);
	s_in2(35,21)            <= s_out2(36,22);
	s_locks_lower_in(35,21) <= s_locks_lower_out(36,21);

		normal_cell_35_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,22),
			fetch              => s_fetch(35,22),
			data_in            => s_data_in(35,22),
			data_out           => s_data_out(35,22),
			out1               => s_out1(35,22),
			out2               => s_out2(35,22),
			lock_lower_row_out => s_locks_lower_out(35,22),
			lock_lower_row_in  => s_locks_lower_in(35,22),
			in1                => s_in1(35,22),
			in2                => s_in2(35,22),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(22)
		);
	s_in1(35,22)            <= s_out1(36,22);
	s_in2(35,22)            <= s_out2(36,23);
	s_locks_lower_in(35,22) <= s_locks_lower_out(36,22);

		normal_cell_35_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,23),
			fetch              => s_fetch(35,23),
			data_in            => s_data_in(35,23),
			data_out           => s_data_out(35,23),
			out1               => s_out1(35,23),
			out2               => s_out2(35,23),
			lock_lower_row_out => s_locks_lower_out(35,23),
			lock_lower_row_in  => s_locks_lower_in(35,23),
			in1                => s_in1(35,23),
			in2                => s_in2(35,23),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(23)
		);
	s_in1(35,23)            <= s_out1(36,23);
	s_in2(35,23)            <= s_out2(36,24);
	s_locks_lower_in(35,23) <= s_locks_lower_out(36,23);

		normal_cell_35_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,24),
			fetch              => s_fetch(35,24),
			data_in            => s_data_in(35,24),
			data_out           => s_data_out(35,24),
			out1               => s_out1(35,24),
			out2               => s_out2(35,24),
			lock_lower_row_out => s_locks_lower_out(35,24),
			lock_lower_row_in  => s_locks_lower_in(35,24),
			in1                => s_in1(35,24),
			in2                => s_in2(35,24),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(24)
		);
	s_in1(35,24)            <= s_out1(36,24);
	s_in2(35,24)            <= s_out2(36,25);
	s_locks_lower_in(35,24) <= s_locks_lower_out(36,24);

		normal_cell_35_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,25),
			fetch              => s_fetch(35,25),
			data_in            => s_data_in(35,25),
			data_out           => s_data_out(35,25),
			out1               => s_out1(35,25),
			out2               => s_out2(35,25),
			lock_lower_row_out => s_locks_lower_out(35,25),
			lock_lower_row_in  => s_locks_lower_in(35,25),
			in1                => s_in1(35,25),
			in2                => s_in2(35,25),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(25)
		);
	s_in1(35,25)            <= s_out1(36,25);
	s_in2(35,25)            <= s_out2(36,26);
	s_locks_lower_in(35,25) <= s_locks_lower_out(36,25);

		normal_cell_35_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,26),
			fetch              => s_fetch(35,26),
			data_in            => s_data_in(35,26),
			data_out           => s_data_out(35,26),
			out1               => s_out1(35,26),
			out2               => s_out2(35,26),
			lock_lower_row_out => s_locks_lower_out(35,26),
			lock_lower_row_in  => s_locks_lower_in(35,26),
			in1                => s_in1(35,26),
			in2                => s_in2(35,26),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(26)
		);
	s_in1(35,26)            <= s_out1(36,26);
	s_in2(35,26)            <= s_out2(36,27);
	s_locks_lower_in(35,26) <= s_locks_lower_out(36,26);

		normal_cell_35_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,27),
			fetch              => s_fetch(35,27),
			data_in            => s_data_in(35,27),
			data_out           => s_data_out(35,27),
			out1               => s_out1(35,27),
			out2               => s_out2(35,27),
			lock_lower_row_out => s_locks_lower_out(35,27),
			lock_lower_row_in  => s_locks_lower_in(35,27),
			in1                => s_in1(35,27),
			in2                => s_in2(35,27),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(27)
		);
	s_in1(35,27)            <= s_out1(36,27);
	s_in2(35,27)            <= s_out2(36,28);
	s_locks_lower_in(35,27) <= s_locks_lower_out(36,27);

		normal_cell_35_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,28),
			fetch              => s_fetch(35,28),
			data_in            => s_data_in(35,28),
			data_out           => s_data_out(35,28),
			out1               => s_out1(35,28),
			out2               => s_out2(35,28),
			lock_lower_row_out => s_locks_lower_out(35,28),
			lock_lower_row_in  => s_locks_lower_in(35,28),
			in1                => s_in1(35,28),
			in2                => s_in2(35,28),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(28)
		);
	s_in1(35,28)            <= s_out1(36,28);
	s_in2(35,28)            <= s_out2(36,29);
	s_locks_lower_in(35,28) <= s_locks_lower_out(36,28);

		normal_cell_35_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,29),
			fetch              => s_fetch(35,29),
			data_in            => s_data_in(35,29),
			data_out           => s_data_out(35,29),
			out1               => s_out1(35,29),
			out2               => s_out2(35,29),
			lock_lower_row_out => s_locks_lower_out(35,29),
			lock_lower_row_in  => s_locks_lower_in(35,29),
			in1                => s_in1(35,29),
			in2                => s_in2(35,29),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(29)
		);
	s_in1(35,29)            <= s_out1(36,29);
	s_in2(35,29)            <= s_out2(36,30);
	s_locks_lower_in(35,29) <= s_locks_lower_out(36,29);

		normal_cell_35_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,30),
			fetch              => s_fetch(35,30),
			data_in            => s_data_in(35,30),
			data_out           => s_data_out(35,30),
			out1               => s_out1(35,30),
			out2               => s_out2(35,30),
			lock_lower_row_out => s_locks_lower_out(35,30),
			lock_lower_row_in  => s_locks_lower_in(35,30),
			in1                => s_in1(35,30),
			in2                => s_in2(35,30),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(30)
		);
	s_in1(35,30)            <= s_out1(36,30);
	s_in2(35,30)            <= s_out2(36,31);
	s_locks_lower_in(35,30) <= s_locks_lower_out(36,30);

		normal_cell_35_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,31),
			fetch              => s_fetch(35,31),
			data_in            => s_data_in(35,31),
			data_out           => s_data_out(35,31),
			out1               => s_out1(35,31),
			out2               => s_out2(35,31),
			lock_lower_row_out => s_locks_lower_out(35,31),
			lock_lower_row_in  => s_locks_lower_in(35,31),
			in1                => s_in1(35,31),
			in2                => s_in2(35,31),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(31)
		);
	s_in1(35,31)            <= s_out1(36,31);
	s_in2(35,31)            <= s_out2(36,32);
	s_locks_lower_in(35,31) <= s_locks_lower_out(36,31);

		normal_cell_35_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,32),
			fetch              => s_fetch(35,32),
			data_in            => s_data_in(35,32),
			data_out           => s_data_out(35,32),
			out1               => s_out1(35,32),
			out2               => s_out2(35,32),
			lock_lower_row_out => s_locks_lower_out(35,32),
			lock_lower_row_in  => s_locks_lower_in(35,32),
			in1                => s_in1(35,32),
			in2                => s_in2(35,32),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(32)
		);
	s_in1(35,32)            <= s_out1(36,32);
	s_in2(35,32)            <= s_out2(36,33);
	s_locks_lower_in(35,32) <= s_locks_lower_out(36,32);

		normal_cell_35_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,33),
			fetch              => s_fetch(35,33),
			data_in            => s_data_in(35,33),
			data_out           => s_data_out(35,33),
			out1               => s_out1(35,33),
			out2               => s_out2(35,33),
			lock_lower_row_out => s_locks_lower_out(35,33),
			lock_lower_row_in  => s_locks_lower_in(35,33),
			in1                => s_in1(35,33),
			in2                => s_in2(35,33),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(33)
		);
	s_in1(35,33)            <= s_out1(36,33);
	s_in2(35,33)            <= s_out2(36,34);
	s_locks_lower_in(35,33) <= s_locks_lower_out(36,33);

		normal_cell_35_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,34),
			fetch              => s_fetch(35,34),
			data_in            => s_data_in(35,34),
			data_out           => s_data_out(35,34),
			out1               => s_out1(35,34),
			out2               => s_out2(35,34),
			lock_lower_row_out => s_locks_lower_out(35,34),
			lock_lower_row_in  => s_locks_lower_in(35,34),
			in1                => s_in1(35,34),
			in2                => s_in2(35,34),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(34)
		);
	s_in1(35,34)            <= s_out1(36,34);
	s_in2(35,34)            <= s_out2(36,35);
	s_locks_lower_in(35,34) <= s_locks_lower_out(36,34);

		normal_cell_35_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,35),
			fetch              => s_fetch(35,35),
			data_in            => s_data_in(35,35),
			data_out           => s_data_out(35,35),
			out1               => s_out1(35,35),
			out2               => s_out2(35,35),
			lock_lower_row_out => s_locks_lower_out(35,35),
			lock_lower_row_in  => s_locks_lower_in(35,35),
			in1                => s_in1(35,35),
			in2                => s_in2(35,35),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(35)
		);
	s_in1(35,35)            <= s_out1(36,35);
	s_in2(35,35)            <= s_out2(36,36);
	s_locks_lower_in(35,35) <= s_locks_lower_out(36,35);

		normal_cell_35_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,36),
			fetch              => s_fetch(35,36),
			data_in            => s_data_in(35,36),
			data_out           => s_data_out(35,36),
			out1               => s_out1(35,36),
			out2               => s_out2(35,36),
			lock_lower_row_out => s_locks_lower_out(35,36),
			lock_lower_row_in  => s_locks_lower_in(35,36),
			in1                => s_in1(35,36),
			in2                => s_in2(35,36),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(36)
		);
	s_in1(35,36)            <= s_out1(36,36);
	s_in2(35,36)            <= s_out2(36,37);
	s_locks_lower_in(35,36) <= s_locks_lower_out(36,36);

		normal_cell_35_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,37),
			fetch              => s_fetch(35,37),
			data_in            => s_data_in(35,37),
			data_out           => s_data_out(35,37),
			out1               => s_out1(35,37),
			out2               => s_out2(35,37),
			lock_lower_row_out => s_locks_lower_out(35,37),
			lock_lower_row_in  => s_locks_lower_in(35,37),
			in1                => s_in1(35,37),
			in2                => s_in2(35,37),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(37)
		);
	s_in1(35,37)            <= s_out1(36,37);
	s_in2(35,37)            <= s_out2(36,38);
	s_locks_lower_in(35,37) <= s_locks_lower_out(36,37);

		normal_cell_35_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,38),
			fetch              => s_fetch(35,38),
			data_in            => s_data_in(35,38),
			data_out           => s_data_out(35,38),
			out1               => s_out1(35,38),
			out2               => s_out2(35,38),
			lock_lower_row_out => s_locks_lower_out(35,38),
			lock_lower_row_in  => s_locks_lower_in(35,38),
			in1                => s_in1(35,38),
			in2                => s_in2(35,38),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(38)
		);
	s_in1(35,38)            <= s_out1(36,38);
	s_in2(35,38)            <= s_out2(36,39);
	s_locks_lower_in(35,38) <= s_locks_lower_out(36,38);

		normal_cell_35_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,39),
			fetch              => s_fetch(35,39),
			data_in            => s_data_in(35,39),
			data_out           => s_data_out(35,39),
			out1               => s_out1(35,39),
			out2               => s_out2(35,39),
			lock_lower_row_out => s_locks_lower_out(35,39),
			lock_lower_row_in  => s_locks_lower_in(35,39),
			in1                => s_in1(35,39),
			in2                => s_in2(35,39),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(39)
		);
	s_in1(35,39)            <= s_out1(36,39);
	s_in2(35,39)            <= s_out2(36,40);
	s_locks_lower_in(35,39) <= s_locks_lower_out(36,39);

		normal_cell_35_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,40),
			fetch              => s_fetch(35,40),
			data_in            => s_data_in(35,40),
			data_out           => s_data_out(35,40),
			out1               => s_out1(35,40),
			out2               => s_out2(35,40),
			lock_lower_row_out => s_locks_lower_out(35,40),
			lock_lower_row_in  => s_locks_lower_in(35,40),
			in1                => s_in1(35,40),
			in2                => s_in2(35,40),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(40)
		);
	s_in1(35,40)            <= s_out1(36,40);
	s_in2(35,40)            <= s_out2(36,41);
	s_locks_lower_in(35,40) <= s_locks_lower_out(36,40);

		normal_cell_35_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,41),
			fetch              => s_fetch(35,41),
			data_in            => s_data_in(35,41),
			data_out           => s_data_out(35,41),
			out1               => s_out1(35,41),
			out2               => s_out2(35,41),
			lock_lower_row_out => s_locks_lower_out(35,41),
			lock_lower_row_in  => s_locks_lower_in(35,41),
			in1                => s_in1(35,41),
			in2                => s_in2(35,41),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(41)
		);
	s_in1(35,41)            <= s_out1(36,41);
	s_in2(35,41)            <= s_out2(36,42);
	s_locks_lower_in(35,41) <= s_locks_lower_out(36,41);

		normal_cell_35_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,42),
			fetch              => s_fetch(35,42),
			data_in            => s_data_in(35,42),
			data_out           => s_data_out(35,42),
			out1               => s_out1(35,42),
			out2               => s_out2(35,42),
			lock_lower_row_out => s_locks_lower_out(35,42),
			lock_lower_row_in  => s_locks_lower_in(35,42),
			in1                => s_in1(35,42),
			in2                => s_in2(35,42),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(42)
		);
	s_in1(35,42)            <= s_out1(36,42);
	s_in2(35,42)            <= s_out2(36,43);
	s_locks_lower_in(35,42) <= s_locks_lower_out(36,42);

		normal_cell_35_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,43),
			fetch              => s_fetch(35,43),
			data_in            => s_data_in(35,43),
			data_out           => s_data_out(35,43),
			out1               => s_out1(35,43),
			out2               => s_out2(35,43),
			lock_lower_row_out => s_locks_lower_out(35,43),
			lock_lower_row_in  => s_locks_lower_in(35,43),
			in1                => s_in1(35,43),
			in2                => s_in2(35,43),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(43)
		);
	s_in1(35,43)            <= s_out1(36,43);
	s_in2(35,43)            <= s_out2(36,44);
	s_locks_lower_in(35,43) <= s_locks_lower_out(36,43);

		normal_cell_35_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,44),
			fetch              => s_fetch(35,44),
			data_in            => s_data_in(35,44),
			data_out           => s_data_out(35,44),
			out1               => s_out1(35,44),
			out2               => s_out2(35,44),
			lock_lower_row_out => s_locks_lower_out(35,44),
			lock_lower_row_in  => s_locks_lower_in(35,44),
			in1                => s_in1(35,44),
			in2                => s_in2(35,44),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(44)
		);
	s_in1(35,44)            <= s_out1(36,44);
	s_in2(35,44)            <= s_out2(36,45);
	s_locks_lower_in(35,44) <= s_locks_lower_out(36,44);

		normal_cell_35_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,45),
			fetch              => s_fetch(35,45),
			data_in            => s_data_in(35,45),
			data_out           => s_data_out(35,45),
			out1               => s_out1(35,45),
			out2               => s_out2(35,45),
			lock_lower_row_out => s_locks_lower_out(35,45),
			lock_lower_row_in  => s_locks_lower_in(35,45),
			in1                => s_in1(35,45),
			in2                => s_in2(35,45),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(45)
		);
	s_in1(35,45)            <= s_out1(36,45);
	s_in2(35,45)            <= s_out2(36,46);
	s_locks_lower_in(35,45) <= s_locks_lower_out(36,45);

		normal_cell_35_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,46),
			fetch              => s_fetch(35,46),
			data_in            => s_data_in(35,46),
			data_out           => s_data_out(35,46),
			out1               => s_out1(35,46),
			out2               => s_out2(35,46),
			lock_lower_row_out => s_locks_lower_out(35,46),
			lock_lower_row_in  => s_locks_lower_in(35,46),
			in1                => s_in1(35,46),
			in2                => s_in2(35,46),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(46)
		);
	s_in1(35,46)            <= s_out1(36,46);
	s_in2(35,46)            <= s_out2(36,47);
	s_locks_lower_in(35,46) <= s_locks_lower_out(36,46);

		normal_cell_35_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,47),
			fetch              => s_fetch(35,47),
			data_in            => s_data_in(35,47),
			data_out           => s_data_out(35,47),
			out1               => s_out1(35,47),
			out2               => s_out2(35,47),
			lock_lower_row_out => s_locks_lower_out(35,47),
			lock_lower_row_in  => s_locks_lower_in(35,47),
			in1                => s_in1(35,47),
			in2                => s_in2(35,47),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(47)
		);
	s_in1(35,47)            <= s_out1(36,47);
	s_in2(35,47)            <= s_out2(36,48);
	s_locks_lower_in(35,47) <= s_locks_lower_out(36,47);

		normal_cell_35_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,48),
			fetch              => s_fetch(35,48),
			data_in            => s_data_in(35,48),
			data_out           => s_data_out(35,48),
			out1               => s_out1(35,48),
			out2               => s_out2(35,48),
			lock_lower_row_out => s_locks_lower_out(35,48),
			lock_lower_row_in  => s_locks_lower_in(35,48),
			in1                => s_in1(35,48),
			in2                => s_in2(35,48),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(48)
		);
	s_in1(35,48)            <= s_out1(36,48);
	s_in2(35,48)            <= s_out2(36,49);
	s_locks_lower_in(35,48) <= s_locks_lower_out(36,48);

		normal_cell_35_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,49),
			fetch              => s_fetch(35,49),
			data_in            => s_data_in(35,49),
			data_out           => s_data_out(35,49),
			out1               => s_out1(35,49),
			out2               => s_out2(35,49),
			lock_lower_row_out => s_locks_lower_out(35,49),
			lock_lower_row_in  => s_locks_lower_in(35,49),
			in1                => s_in1(35,49),
			in2                => s_in2(35,49),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(49)
		);
	s_in1(35,49)            <= s_out1(36,49);
	s_in2(35,49)            <= s_out2(36,50);
	s_locks_lower_in(35,49) <= s_locks_lower_out(36,49);

		normal_cell_35_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,50),
			fetch              => s_fetch(35,50),
			data_in            => s_data_in(35,50),
			data_out           => s_data_out(35,50),
			out1               => s_out1(35,50),
			out2               => s_out2(35,50),
			lock_lower_row_out => s_locks_lower_out(35,50),
			lock_lower_row_in  => s_locks_lower_in(35,50),
			in1                => s_in1(35,50),
			in2                => s_in2(35,50),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(50)
		);
	s_in1(35,50)            <= s_out1(36,50);
	s_in2(35,50)            <= s_out2(36,51);
	s_locks_lower_in(35,50) <= s_locks_lower_out(36,50);

		normal_cell_35_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,51),
			fetch              => s_fetch(35,51),
			data_in            => s_data_in(35,51),
			data_out           => s_data_out(35,51),
			out1               => s_out1(35,51),
			out2               => s_out2(35,51),
			lock_lower_row_out => s_locks_lower_out(35,51),
			lock_lower_row_in  => s_locks_lower_in(35,51),
			in1                => s_in1(35,51),
			in2                => s_in2(35,51),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(51)
		);
	s_in1(35,51)            <= s_out1(36,51);
	s_in2(35,51)            <= s_out2(36,52);
	s_locks_lower_in(35,51) <= s_locks_lower_out(36,51);

		normal_cell_35_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,52),
			fetch              => s_fetch(35,52),
			data_in            => s_data_in(35,52),
			data_out           => s_data_out(35,52),
			out1               => s_out1(35,52),
			out2               => s_out2(35,52),
			lock_lower_row_out => s_locks_lower_out(35,52),
			lock_lower_row_in  => s_locks_lower_in(35,52),
			in1                => s_in1(35,52),
			in2                => s_in2(35,52),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(52)
		);
	s_in1(35,52)            <= s_out1(36,52);
	s_in2(35,52)            <= s_out2(36,53);
	s_locks_lower_in(35,52) <= s_locks_lower_out(36,52);

		normal_cell_35_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,53),
			fetch              => s_fetch(35,53),
			data_in            => s_data_in(35,53),
			data_out           => s_data_out(35,53),
			out1               => s_out1(35,53),
			out2               => s_out2(35,53),
			lock_lower_row_out => s_locks_lower_out(35,53),
			lock_lower_row_in  => s_locks_lower_in(35,53),
			in1                => s_in1(35,53),
			in2                => s_in2(35,53),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(53)
		);
	s_in1(35,53)            <= s_out1(36,53);
	s_in2(35,53)            <= s_out2(36,54);
	s_locks_lower_in(35,53) <= s_locks_lower_out(36,53);

		normal_cell_35_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,54),
			fetch              => s_fetch(35,54),
			data_in            => s_data_in(35,54),
			data_out           => s_data_out(35,54),
			out1               => s_out1(35,54),
			out2               => s_out2(35,54),
			lock_lower_row_out => s_locks_lower_out(35,54),
			lock_lower_row_in  => s_locks_lower_in(35,54),
			in1                => s_in1(35,54),
			in2                => s_in2(35,54),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(54)
		);
	s_in1(35,54)            <= s_out1(36,54);
	s_in2(35,54)            <= s_out2(36,55);
	s_locks_lower_in(35,54) <= s_locks_lower_out(36,54);

		normal_cell_35_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,55),
			fetch              => s_fetch(35,55),
			data_in            => s_data_in(35,55),
			data_out           => s_data_out(35,55),
			out1               => s_out1(35,55),
			out2               => s_out2(35,55),
			lock_lower_row_out => s_locks_lower_out(35,55),
			lock_lower_row_in  => s_locks_lower_in(35,55),
			in1                => s_in1(35,55),
			in2                => s_in2(35,55),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(55)
		);
	s_in1(35,55)            <= s_out1(36,55);
	s_in2(35,55)            <= s_out2(36,56);
	s_locks_lower_in(35,55) <= s_locks_lower_out(36,55);

		normal_cell_35_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,56),
			fetch              => s_fetch(35,56),
			data_in            => s_data_in(35,56),
			data_out           => s_data_out(35,56),
			out1               => s_out1(35,56),
			out2               => s_out2(35,56),
			lock_lower_row_out => s_locks_lower_out(35,56),
			lock_lower_row_in  => s_locks_lower_in(35,56),
			in1                => s_in1(35,56),
			in2                => s_in2(35,56),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(56)
		);
	s_in1(35,56)            <= s_out1(36,56);
	s_in2(35,56)            <= s_out2(36,57);
	s_locks_lower_in(35,56) <= s_locks_lower_out(36,56);

		normal_cell_35_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,57),
			fetch              => s_fetch(35,57),
			data_in            => s_data_in(35,57),
			data_out           => s_data_out(35,57),
			out1               => s_out1(35,57),
			out2               => s_out2(35,57),
			lock_lower_row_out => s_locks_lower_out(35,57),
			lock_lower_row_in  => s_locks_lower_in(35,57),
			in1                => s_in1(35,57),
			in2                => s_in2(35,57),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(57)
		);
	s_in1(35,57)            <= s_out1(36,57);
	s_in2(35,57)            <= s_out2(36,58);
	s_locks_lower_in(35,57) <= s_locks_lower_out(36,57);

		normal_cell_35_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,58),
			fetch              => s_fetch(35,58),
			data_in            => s_data_in(35,58),
			data_out           => s_data_out(35,58),
			out1               => s_out1(35,58),
			out2               => s_out2(35,58),
			lock_lower_row_out => s_locks_lower_out(35,58),
			lock_lower_row_in  => s_locks_lower_in(35,58),
			in1                => s_in1(35,58),
			in2                => s_in2(35,58),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(58)
		);
	s_in1(35,58)            <= s_out1(36,58);
	s_in2(35,58)            <= s_out2(36,59);
	s_locks_lower_in(35,58) <= s_locks_lower_out(36,58);

		normal_cell_35_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,59),
			fetch              => s_fetch(35,59),
			data_in            => s_data_in(35,59),
			data_out           => s_data_out(35,59),
			out1               => s_out1(35,59),
			out2               => s_out2(35,59),
			lock_lower_row_out => s_locks_lower_out(35,59),
			lock_lower_row_in  => s_locks_lower_in(35,59),
			in1                => s_in1(35,59),
			in2                => s_in2(35,59),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(59)
		);
	s_in1(35,59)            <= s_out1(36,59);
	s_in2(35,59)            <= s_out2(36,60);
	s_locks_lower_in(35,59) <= s_locks_lower_out(36,59);

		last_col_cell_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(35,60),
			fetch              => s_fetch(35,60),
			data_in            => s_data_in(35,60),
			data_out           => s_data_out(35,60),
			out1               => s_out1(35,60),
			out2               => s_out2(35,60),
			lock_lower_row_out => s_locks_lower_out(35,60),
			lock_lower_row_in  => s_locks_lower_in(35,60),
			in1                => s_in1(35,60),
			in2                => (others => '0'),
			lock_row           => s_locks(35),
			piv_found          => s_piv_found,
			row_data           => s_row_data(35),
			col_data           => s_col_data(60)
		);
	s_in1(35,60)            <= s_out1(36,60);
	s_locks_lower_in(35,60) <= s_locks_lower_out(36,60);

		normal_cell_36_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,1),
			fetch              => s_fetch(36,1),
			data_in            => s_data_in(36,1),
			data_out           => s_data_out(36,1),
			out1               => s_out1(36,1),
			out2               => s_out2(36,1),
			lock_lower_row_out => s_locks_lower_out(36,1),
			lock_lower_row_in  => s_locks_lower_in(36,1),
			in1                => s_in1(36,1),
			in2                => s_in2(36,1),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(1)
		);
	s_in1(36,1)            <= s_out1(37,1);
	s_in2(36,1)            <= s_out2(37,2);
	s_locks_lower_in(36,1) <= s_locks_lower_out(37,1);

		normal_cell_36_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,2),
			fetch              => s_fetch(36,2),
			data_in            => s_data_in(36,2),
			data_out           => s_data_out(36,2),
			out1               => s_out1(36,2),
			out2               => s_out2(36,2),
			lock_lower_row_out => s_locks_lower_out(36,2),
			lock_lower_row_in  => s_locks_lower_in(36,2),
			in1                => s_in1(36,2),
			in2                => s_in2(36,2),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(2)
		);
	s_in1(36,2)            <= s_out1(37,2);
	s_in2(36,2)            <= s_out2(37,3);
	s_locks_lower_in(36,2) <= s_locks_lower_out(37,2);

		normal_cell_36_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,3),
			fetch              => s_fetch(36,3),
			data_in            => s_data_in(36,3),
			data_out           => s_data_out(36,3),
			out1               => s_out1(36,3),
			out2               => s_out2(36,3),
			lock_lower_row_out => s_locks_lower_out(36,3),
			lock_lower_row_in  => s_locks_lower_in(36,3),
			in1                => s_in1(36,3),
			in2                => s_in2(36,3),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(3)
		);
	s_in1(36,3)            <= s_out1(37,3);
	s_in2(36,3)            <= s_out2(37,4);
	s_locks_lower_in(36,3) <= s_locks_lower_out(37,3);

		normal_cell_36_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,4),
			fetch              => s_fetch(36,4),
			data_in            => s_data_in(36,4),
			data_out           => s_data_out(36,4),
			out1               => s_out1(36,4),
			out2               => s_out2(36,4),
			lock_lower_row_out => s_locks_lower_out(36,4),
			lock_lower_row_in  => s_locks_lower_in(36,4),
			in1                => s_in1(36,4),
			in2                => s_in2(36,4),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(4)
		);
	s_in1(36,4)            <= s_out1(37,4);
	s_in2(36,4)            <= s_out2(37,5);
	s_locks_lower_in(36,4) <= s_locks_lower_out(37,4);

		normal_cell_36_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,5),
			fetch              => s_fetch(36,5),
			data_in            => s_data_in(36,5),
			data_out           => s_data_out(36,5),
			out1               => s_out1(36,5),
			out2               => s_out2(36,5),
			lock_lower_row_out => s_locks_lower_out(36,5),
			lock_lower_row_in  => s_locks_lower_in(36,5),
			in1                => s_in1(36,5),
			in2                => s_in2(36,5),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(5)
		);
	s_in1(36,5)            <= s_out1(37,5);
	s_in2(36,5)            <= s_out2(37,6);
	s_locks_lower_in(36,5) <= s_locks_lower_out(37,5);

		normal_cell_36_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,6),
			fetch              => s_fetch(36,6),
			data_in            => s_data_in(36,6),
			data_out           => s_data_out(36,6),
			out1               => s_out1(36,6),
			out2               => s_out2(36,6),
			lock_lower_row_out => s_locks_lower_out(36,6),
			lock_lower_row_in  => s_locks_lower_in(36,6),
			in1                => s_in1(36,6),
			in2                => s_in2(36,6),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(6)
		);
	s_in1(36,6)            <= s_out1(37,6);
	s_in2(36,6)            <= s_out2(37,7);
	s_locks_lower_in(36,6) <= s_locks_lower_out(37,6);

		normal_cell_36_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,7),
			fetch              => s_fetch(36,7),
			data_in            => s_data_in(36,7),
			data_out           => s_data_out(36,7),
			out1               => s_out1(36,7),
			out2               => s_out2(36,7),
			lock_lower_row_out => s_locks_lower_out(36,7),
			lock_lower_row_in  => s_locks_lower_in(36,7),
			in1                => s_in1(36,7),
			in2                => s_in2(36,7),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(7)
		);
	s_in1(36,7)            <= s_out1(37,7);
	s_in2(36,7)            <= s_out2(37,8);
	s_locks_lower_in(36,7) <= s_locks_lower_out(37,7);

		normal_cell_36_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,8),
			fetch              => s_fetch(36,8),
			data_in            => s_data_in(36,8),
			data_out           => s_data_out(36,8),
			out1               => s_out1(36,8),
			out2               => s_out2(36,8),
			lock_lower_row_out => s_locks_lower_out(36,8),
			lock_lower_row_in  => s_locks_lower_in(36,8),
			in1                => s_in1(36,8),
			in2                => s_in2(36,8),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(8)
		);
	s_in1(36,8)            <= s_out1(37,8);
	s_in2(36,8)            <= s_out2(37,9);
	s_locks_lower_in(36,8) <= s_locks_lower_out(37,8);

		normal_cell_36_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,9),
			fetch              => s_fetch(36,9),
			data_in            => s_data_in(36,9),
			data_out           => s_data_out(36,9),
			out1               => s_out1(36,9),
			out2               => s_out2(36,9),
			lock_lower_row_out => s_locks_lower_out(36,9),
			lock_lower_row_in  => s_locks_lower_in(36,9),
			in1                => s_in1(36,9),
			in2                => s_in2(36,9),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(9)
		);
	s_in1(36,9)            <= s_out1(37,9);
	s_in2(36,9)            <= s_out2(37,10);
	s_locks_lower_in(36,9) <= s_locks_lower_out(37,9);

		normal_cell_36_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,10),
			fetch              => s_fetch(36,10),
			data_in            => s_data_in(36,10),
			data_out           => s_data_out(36,10),
			out1               => s_out1(36,10),
			out2               => s_out2(36,10),
			lock_lower_row_out => s_locks_lower_out(36,10),
			lock_lower_row_in  => s_locks_lower_in(36,10),
			in1                => s_in1(36,10),
			in2                => s_in2(36,10),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(10)
		);
	s_in1(36,10)            <= s_out1(37,10);
	s_in2(36,10)            <= s_out2(37,11);
	s_locks_lower_in(36,10) <= s_locks_lower_out(37,10);

		normal_cell_36_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,11),
			fetch              => s_fetch(36,11),
			data_in            => s_data_in(36,11),
			data_out           => s_data_out(36,11),
			out1               => s_out1(36,11),
			out2               => s_out2(36,11),
			lock_lower_row_out => s_locks_lower_out(36,11),
			lock_lower_row_in  => s_locks_lower_in(36,11),
			in1                => s_in1(36,11),
			in2                => s_in2(36,11),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(11)
		);
	s_in1(36,11)            <= s_out1(37,11);
	s_in2(36,11)            <= s_out2(37,12);
	s_locks_lower_in(36,11) <= s_locks_lower_out(37,11);

		normal_cell_36_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,12),
			fetch              => s_fetch(36,12),
			data_in            => s_data_in(36,12),
			data_out           => s_data_out(36,12),
			out1               => s_out1(36,12),
			out2               => s_out2(36,12),
			lock_lower_row_out => s_locks_lower_out(36,12),
			lock_lower_row_in  => s_locks_lower_in(36,12),
			in1                => s_in1(36,12),
			in2                => s_in2(36,12),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(12)
		);
	s_in1(36,12)            <= s_out1(37,12);
	s_in2(36,12)            <= s_out2(37,13);
	s_locks_lower_in(36,12) <= s_locks_lower_out(37,12);

		normal_cell_36_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,13),
			fetch              => s_fetch(36,13),
			data_in            => s_data_in(36,13),
			data_out           => s_data_out(36,13),
			out1               => s_out1(36,13),
			out2               => s_out2(36,13),
			lock_lower_row_out => s_locks_lower_out(36,13),
			lock_lower_row_in  => s_locks_lower_in(36,13),
			in1                => s_in1(36,13),
			in2                => s_in2(36,13),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(13)
		);
	s_in1(36,13)            <= s_out1(37,13);
	s_in2(36,13)            <= s_out2(37,14);
	s_locks_lower_in(36,13) <= s_locks_lower_out(37,13);

		normal_cell_36_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,14),
			fetch              => s_fetch(36,14),
			data_in            => s_data_in(36,14),
			data_out           => s_data_out(36,14),
			out1               => s_out1(36,14),
			out2               => s_out2(36,14),
			lock_lower_row_out => s_locks_lower_out(36,14),
			lock_lower_row_in  => s_locks_lower_in(36,14),
			in1                => s_in1(36,14),
			in2                => s_in2(36,14),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(14)
		);
	s_in1(36,14)            <= s_out1(37,14);
	s_in2(36,14)            <= s_out2(37,15);
	s_locks_lower_in(36,14) <= s_locks_lower_out(37,14);

		normal_cell_36_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,15),
			fetch              => s_fetch(36,15),
			data_in            => s_data_in(36,15),
			data_out           => s_data_out(36,15),
			out1               => s_out1(36,15),
			out2               => s_out2(36,15),
			lock_lower_row_out => s_locks_lower_out(36,15),
			lock_lower_row_in  => s_locks_lower_in(36,15),
			in1                => s_in1(36,15),
			in2                => s_in2(36,15),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(15)
		);
	s_in1(36,15)            <= s_out1(37,15);
	s_in2(36,15)            <= s_out2(37,16);
	s_locks_lower_in(36,15) <= s_locks_lower_out(37,15);

		normal_cell_36_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,16),
			fetch              => s_fetch(36,16),
			data_in            => s_data_in(36,16),
			data_out           => s_data_out(36,16),
			out1               => s_out1(36,16),
			out2               => s_out2(36,16),
			lock_lower_row_out => s_locks_lower_out(36,16),
			lock_lower_row_in  => s_locks_lower_in(36,16),
			in1                => s_in1(36,16),
			in2                => s_in2(36,16),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(16)
		);
	s_in1(36,16)            <= s_out1(37,16);
	s_in2(36,16)            <= s_out2(37,17);
	s_locks_lower_in(36,16) <= s_locks_lower_out(37,16);

		normal_cell_36_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,17),
			fetch              => s_fetch(36,17),
			data_in            => s_data_in(36,17),
			data_out           => s_data_out(36,17),
			out1               => s_out1(36,17),
			out2               => s_out2(36,17),
			lock_lower_row_out => s_locks_lower_out(36,17),
			lock_lower_row_in  => s_locks_lower_in(36,17),
			in1                => s_in1(36,17),
			in2                => s_in2(36,17),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(17)
		);
	s_in1(36,17)            <= s_out1(37,17);
	s_in2(36,17)            <= s_out2(37,18);
	s_locks_lower_in(36,17) <= s_locks_lower_out(37,17);

		normal_cell_36_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,18),
			fetch              => s_fetch(36,18),
			data_in            => s_data_in(36,18),
			data_out           => s_data_out(36,18),
			out1               => s_out1(36,18),
			out2               => s_out2(36,18),
			lock_lower_row_out => s_locks_lower_out(36,18),
			lock_lower_row_in  => s_locks_lower_in(36,18),
			in1                => s_in1(36,18),
			in2                => s_in2(36,18),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(18)
		);
	s_in1(36,18)            <= s_out1(37,18);
	s_in2(36,18)            <= s_out2(37,19);
	s_locks_lower_in(36,18) <= s_locks_lower_out(37,18);

		normal_cell_36_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,19),
			fetch              => s_fetch(36,19),
			data_in            => s_data_in(36,19),
			data_out           => s_data_out(36,19),
			out1               => s_out1(36,19),
			out2               => s_out2(36,19),
			lock_lower_row_out => s_locks_lower_out(36,19),
			lock_lower_row_in  => s_locks_lower_in(36,19),
			in1                => s_in1(36,19),
			in2                => s_in2(36,19),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(19)
		);
	s_in1(36,19)            <= s_out1(37,19);
	s_in2(36,19)            <= s_out2(37,20);
	s_locks_lower_in(36,19) <= s_locks_lower_out(37,19);

		normal_cell_36_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,20),
			fetch              => s_fetch(36,20),
			data_in            => s_data_in(36,20),
			data_out           => s_data_out(36,20),
			out1               => s_out1(36,20),
			out2               => s_out2(36,20),
			lock_lower_row_out => s_locks_lower_out(36,20),
			lock_lower_row_in  => s_locks_lower_in(36,20),
			in1                => s_in1(36,20),
			in2                => s_in2(36,20),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(20)
		);
	s_in1(36,20)            <= s_out1(37,20);
	s_in2(36,20)            <= s_out2(37,21);
	s_locks_lower_in(36,20) <= s_locks_lower_out(37,20);

		normal_cell_36_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,21),
			fetch              => s_fetch(36,21),
			data_in            => s_data_in(36,21),
			data_out           => s_data_out(36,21),
			out1               => s_out1(36,21),
			out2               => s_out2(36,21),
			lock_lower_row_out => s_locks_lower_out(36,21),
			lock_lower_row_in  => s_locks_lower_in(36,21),
			in1                => s_in1(36,21),
			in2                => s_in2(36,21),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(21)
		);
	s_in1(36,21)            <= s_out1(37,21);
	s_in2(36,21)            <= s_out2(37,22);
	s_locks_lower_in(36,21) <= s_locks_lower_out(37,21);

		normal_cell_36_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,22),
			fetch              => s_fetch(36,22),
			data_in            => s_data_in(36,22),
			data_out           => s_data_out(36,22),
			out1               => s_out1(36,22),
			out2               => s_out2(36,22),
			lock_lower_row_out => s_locks_lower_out(36,22),
			lock_lower_row_in  => s_locks_lower_in(36,22),
			in1                => s_in1(36,22),
			in2                => s_in2(36,22),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(22)
		);
	s_in1(36,22)            <= s_out1(37,22);
	s_in2(36,22)            <= s_out2(37,23);
	s_locks_lower_in(36,22) <= s_locks_lower_out(37,22);

		normal_cell_36_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,23),
			fetch              => s_fetch(36,23),
			data_in            => s_data_in(36,23),
			data_out           => s_data_out(36,23),
			out1               => s_out1(36,23),
			out2               => s_out2(36,23),
			lock_lower_row_out => s_locks_lower_out(36,23),
			lock_lower_row_in  => s_locks_lower_in(36,23),
			in1                => s_in1(36,23),
			in2                => s_in2(36,23),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(23)
		);
	s_in1(36,23)            <= s_out1(37,23);
	s_in2(36,23)            <= s_out2(37,24);
	s_locks_lower_in(36,23) <= s_locks_lower_out(37,23);

		normal_cell_36_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,24),
			fetch              => s_fetch(36,24),
			data_in            => s_data_in(36,24),
			data_out           => s_data_out(36,24),
			out1               => s_out1(36,24),
			out2               => s_out2(36,24),
			lock_lower_row_out => s_locks_lower_out(36,24),
			lock_lower_row_in  => s_locks_lower_in(36,24),
			in1                => s_in1(36,24),
			in2                => s_in2(36,24),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(24)
		);
	s_in1(36,24)            <= s_out1(37,24);
	s_in2(36,24)            <= s_out2(37,25);
	s_locks_lower_in(36,24) <= s_locks_lower_out(37,24);

		normal_cell_36_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,25),
			fetch              => s_fetch(36,25),
			data_in            => s_data_in(36,25),
			data_out           => s_data_out(36,25),
			out1               => s_out1(36,25),
			out2               => s_out2(36,25),
			lock_lower_row_out => s_locks_lower_out(36,25),
			lock_lower_row_in  => s_locks_lower_in(36,25),
			in1                => s_in1(36,25),
			in2                => s_in2(36,25),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(25)
		);
	s_in1(36,25)            <= s_out1(37,25);
	s_in2(36,25)            <= s_out2(37,26);
	s_locks_lower_in(36,25) <= s_locks_lower_out(37,25);

		normal_cell_36_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,26),
			fetch              => s_fetch(36,26),
			data_in            => s_data_in(36,26),
			data_out           => s_data_out(36,26),
			out1               => s_out1(36,26),
			out2               => s_out2(36,26),
			lock_lower_row_out => s_locks_lower_out(36,26),
			lock_lower_row_in  => s_locks_lower_in(36,26),
			in1                => s_in1(36,26),
			in2                => s_in2(36,26),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(26)
		);
	s_in1(36,26)            <= s_out1(37,26);
	s_in2(36,26)            <= s_out2(37,27);
	s_locks_lower_in(36,26) <= s_locks_lower_out(37,26);

		normal_cell_36_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,27),
			fetch              => s_fetch(36,27),
			data_in            => s_data_in(36,27),
			data_out           => s_data_out(36,27),
			out1               => s_out1(36,27),
			out2               => s_out2(36,27),
			lock_lower_row_out => s_locks_lower_out(36,27),
			lock_lower_row_in  => s_locks_lower_in(36,27),
			in1                => s_in1(36,27),
			in2                => s_in2(36,27),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(27)
		);
	s_in1(36,27)            <= s_out1(37,27);
	s_in2(36,27)            <= s_out2(37,28);
	s_locks_lower_in(36,27) <= s_locks_lower_out(37,27);

		normal_cell_36_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,28),
			fetch              => s_fetch(36,28),
			data_in            => s_data_in(36,28),
			data_out           => s_data_out(36,28),
			out1               => s_out1(36,28),
			out2               => s_out2(36,28),
			lock_lower_row_out => s_locks_lower_out(36,28),
			lock_lower_row_in  => s_locks_lower_in(36,28),
			in1                => s_in1(36,28),
			in2                => s_in2(36,28),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(28)
		);
	s_in1(36,28)            <= s_out1(37,28);
	s_in2(36,28)            <= s_out2(37,29);
	s_locks_lower_in(36,28) <= s_locks_lower_out(37,28);

		normal_cell_36_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,29),
			fetch              => s_fetch(36,29),
			data_in            => s_data_in(36,29),
			data_out           => s_data_out(36,29),
			out1               => s_out1(36,29),
			out2               => s_out2(36,29),
			lock_lower_row_out => s_locks_lower_out(36,29),
			lock_lower_row_in  => s_locks_lower_in(36,29),
			in1                => s_in1(36,29),
			in2                => s_in2(36,29),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(29)
		);
	s_in1(36,29)            <= s_out1(37,29);
	s_in2(36,29)            <= s_out2(37,30);
	s_locks_lower_in(36,29) <= s_locks_lower_out(37,29);

		normal_cell_36_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,30),
			fetch              => s_fetch(36,30),
			data_in            => s_data_in(36,30),
			data_out           => s_data_out(36,30),
			out1               => s_out1(36,30),
			out2               => s_out2(36,30),
			lock_lower_row_out => s_locks_lower_out(36,30),
			lock_lower_row_in  => s_locks_lower_in(36,30),
			in1                => s_in1(36,30),
			in2                => s_in2(36,30),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(30)
		);
	s_in1(36,30)            <= s_out1(37,30);
	s_in2(36,30)            <= s_out2(37,31);
	s_locks_lower_in(36,30) <= s_locks_lower_out(37,30);

		normal_cell_36_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,31),
			fetch              => s_fetch(36,31),
			data_in            => s_data_in(36,31),
			data_out           => s_data_out(36,31),
			out1               => s_out1(36,31),
			out2               => s_out2(36,31),
			lock_lower_row_out => s_locks_lower_out(36,31),
			lock_lower_row_in  => s_locks_lower_in(36,31),
			in1                => s_in1(36,31),
			in2                => s_in2(36,31),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(31)
		);
	s_in1(36,31)            <= s_out1(37,31);
	s_in2(36,31)            <= s_out2(37,32);
	s_locks_lower_in(36,31) <= s_locks_lower_out(37,31);

		normal_cell_36_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,32),
			fetch              => s_fetch(36,32),
			data_in            => s_data_in(36,32),
			data_out           => s_data_out(36,32),
			out1               => s_out1(36,32),
			out2               => s_out2(36,32),
			lock_lower_row_out => s_locks_lower_out(36,32),
			lock_lower_row_in  => s_locks_lower_in(36,32),
			in1                => s_in1(36,32),
			in2                => s_in2(36,32),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(32)
		);
	s_in1(36,32)            <= s_out1(37,32);
	s_in2(36,32)            <= s_out2(37,33);
	s_locks_lower_in(36,32) <= s_locks_lower_out(37,32);

		normal_cell_36_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,33),
			fetch              => s_fetch(36,33),
			data_in            => s_data_in(36,33),
			data_out           => s_data_out(36,33),
			out1               => s_out1(36,33),
			out2               => s_out2(36,33),
			lock_lower_row_out => s_locks_lower_out(36,33),
			lock_lower_row_in  => s_locks_lower_in(36,33),
			in1                => s_in1(36,33),
			in2                => s_in2(36,33),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(33)
		);
	s_in1(36,33)            <= s_out1(37,33);
	s_in2(36,33)            <= s_out2(37,34);
	s_locks_lower_in(36,33) <= s_locks_lower_out(37,33);

		normal_cell_36_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,34),
			fetch              => s_fetch(36,34),
			data_in            => s_data_in(36,34),
			data_out           => s_data_out(36,34),
			out1               => s_out1(36,34),
			out2               => s_out2(36,34),
			lock_lower_row_out => s_locks_lower_out(36,34),
			lock_lower_row_in  => s_locks_lower_in(36,34),
			in1                => s_in1(36,34),
			in2                => s_in2(36,34),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(34)
		);
	s_in1(36,34)            <= s_out1(37,34);
	s_in2(36,34)            <= s_out2(37,35);
	s_locks_lower_in(36,34) <= s_locks_lower_out(37,34);

		normal_cell_36_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,35),
			fetch              => s_fetch(36,35),
			data_in            => s_data_in(36,35),
			data_out           => s_data_out(36,35),
			out1               => s_out1(36,35),
			out2               => s_out2(36,35),
			lock_lower_row_out => s_locks_lower_out(36,35),
			lock_lower_row_in  => s_locks_lower_in(36,35),
			in1                => s_in1(36,35),
			in2                => s_in2(36,35),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(35)
		);
	s_in1(36,35)            <= s_out1(37,35);
	s_in2(36,35)            <= s_out2(37,36);
	s_locks_lower_in(36,35) <= s_locks_lower_out(37,35);

		normal_cell_36_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,36),
			fetch              => s_fetch(36,36),
			data_in            => s_data_in(36,36),
			data_out           => s_data_out(36,36),
			out1               => s_out1(36,36),
			out2               => s_out2(36,36),
			lock_lower_row_out => s_locks_lower_out(36,36),
			lock_lower_row_in  => s_locks_lower_in(36,36),
			in1                => s_in1(36,36),
			in2                => s_in2(36,36),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(36)
		);
	s_in1(36,36)            <= s_out1(37,36);
	s_in2(36,36)            <= s_out2(37,37);
	s_locks_lower_in(36,36) <= s_locks_lower_out(37,36);

		normal_cell_36_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,37),
			fetch              => s_fetch(36,37),
			data_in            => s_data_in(36,37),
			data_out           => s_data_out(36,37),
			out1               => s_out1(36,37),
			out2               => s_out2(36,37),
			lock_lower_row_out => s_locks_lower_out(36,37),
			lock_lower_row_in  => s_locks_lower_in(36,37),
			in1                => s_in1(36,37),
			in2                => s_in2(36,37),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(37)
		);
	s_in1(36,37)            <= s_out1(37,37);
	s_in2(36,37)            <= s_out2(37,38);
	s_locks_lower_in(36,37) <= s_locks_lower_out(37,37);

		normal_cell_36_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,38),
			fetch              => s_fetch(36,38),
			data_in            => s_data_in(36,38),
			data_out           => s_data_out(36,38),
			out1               => s_out1(36,38),
			out2               => s_out2(36,38),
			lock_lower_row_out => s_locks_lower_out(36,38),
			lock_lower_row_in  => s_locks_lower_in(36,38),
			in1                => s_in1(36,38),
			in2                => s_in2(36,38),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(38)
		);
	s_in1(36,38)            <= s_out1(37,38);
	s_in2(36,38)            <= s_out2(37,39);
	s_locks_lower_in(36,38) <= s_locks_lower_out(37,38);

		normal_cell_36_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,39),
			fetch              => s_fetch(36,39),
			data_in            => s_data_in(36,39),
			data_out           => s_data_out(36,39),
			out1               => s_out1(36,39),
			out2               => s_out2(36,39),
			lock_lower_row_out => s_locks_lower_out(36,39),
			lock_lower_row_in  => s_locks_lower_in(36,39),
			in1                => s_in1(36,39),
			in2                => s_in2(36,39),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(39)
		);
	s_in1(36,39)            <= s_out1(37,39);
	s_in2(36,39)            <= s_out2(37,40);
	s_locks_lower_in(36,39) <= s_locks_lower_out(37,39);

		normal_cell_36_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,40),
			fetch              => s_fetch(36,40),
			data_in            => s_data_in(36,40),
			data_out           => s_data_out(36,40),
			out1               => s_out1(36,40),
			out2               => s_out2(36,40),
			lock_lower_row_out => s_locks_lower_out(36,40),
			lock_lower_row_in  => s_locks_lower_in(36,40),
			in1                => s_in1(36,40),
			in2                => s_in2(36,40),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(40)
		);
	s_in1(36,40)            <= s_out1(37,40);
	s_in2(36,40)            <= s_out2(37,41);
	s_locks_lower_in(36,40) <= s_locks_lower_out(37,40);

		normal_cell_36_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,41),
			fetch              => s_fetch(36,41),
			data_in            => s_data_in(36,41),
			data_out           => s_data_out(36,41),
			out1               => s_out1(36,41),
			out2               => s_out2(36,41),
			lock_lower_row_out => s_locks_lower_out(36,41),
			lock_lower_row_in  => s_locks_lower_in(36,41),
			in1                => s_in1(36,41),
			in2                => s_in2(36,41),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(41)
		);
	s_in1(36,41)            <= s_out1(37,41);
	s_in2(36,41)            <= s_out2(37,42);
	s_locks_lower_in(36,41) <= s_locks_lower_out(37,41);

		normal_cell_36_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,42),
			fetch              => s_fetch(36,42),
			data_in            => s_data_in(36,42),
			data_out           => s_data_out(36,42),
			out1               => s_out1(36,42),
			out2               => s_out2(36,42),
			lock_lower_row_out => s_locks_lower_out(36,42),
			lock_lower_row_in  => s_locks_lower_in(36,42),
			in1                => s_in1(36,42),
			in2                => s_in2(36,42),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(42)
		);
	s_in1(36,42)            <= s_out1(37,42);
	s_in2(36,42)            <= s_out2(37,43);
	s_locks_lower_in(36,42) <= s_locks_lower_out(37,42);

		normal_cell_36_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,43),
			fetch              => s_fetch(36,43),
			data_in            => s_data_in(36,43),
			data_out           => s_data_out(36,43),
			out1               => s_out1(36,43),
			out2               => s_out2(36,43),
			lock_lower_row_out => s_locks_lower_out(36,43),
			lock_lower_row_in  => s_locks_lower_in(36,43),
			in1                => s_in1(36,43),
			in2                => s_in2(36,43),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(43)
		);
	s_in1(36,43)            <= s_out1(37,43);
	s_in2(36,43)            <= s_out2(37,44);
	s_locks_lower_in(36,43) <= s_locks_lower_out(37,43);

		normal_cell_36_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,44),
			fetch              => s_fetch(36,44),
			data_in            => s_data_in(36,44),
			data_out           => s_data_out(36,44),
			out1               => s_out1(36,44),
			out2               => s_out2(36,44),
			lock_lower_row_out => s_locks_lower_out(36,44),
			lock_lower_row_in  => s_locks_lower_in(36,44),
			in1                => s_in1(36,44),
			in2                => s_in2(36,44),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(44)
		);
	s_in1(36,44)            <= s_out1(37,44);
	s_in2(36,44)            <= s_out2(37,45);
	s_locks_lower_in(36,44) <= s_locks_lower_out(37,44);

		normal_cell_36_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,45),
			fetch              => s_fetch(36,45),
			data_in            => s_data_in(36,45),
			data_out           => s_data_out(36,45),
			out1               => s_out1(36,45),
			out2               => s_out2(36,45),
			lock_lower_row_out => s_locks_lower_out(36,45),
			lock_lower_row_in  => s_locks_lower_in(36,45),
			in1                => s_in1(36,45),
			in2                => s_in2(36,45),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(45)
		);
	s_in1(36,45)            <= s_out1(37,45);
	s_in2(36,45)            <= s_out2(37,46);
	s_locks_lower_in(36,45) <= s_locks_lower_out(37,45);

		normal_cell_36_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,46),
			fetch              => s_fetch(36,46),
			data_in            => s_data_in(36,46),
			data_out           => s_data_out(36,46),
			out1               => s_out1(36,46),
			out2               => s_out2(36,46),
			lock_lower_row_out => s_locks_lower_out(36,46),
			lock_lower_row_in  => s_locks_lower_in(36,46),
			in1                => s_in1(36,46),
			in2                => s_in2(36,46),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(46)
		);
	s_in1(36,46)            <= s_out1(37,46);
	s_in2(36,46)            <= s_out2(37,47);
	s_locks_lower_in(36,46) <= s_locks_lower_out(37,46);

		normal_cell_36_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,47),
			fetch              => s_fetch(36,47),
			data_in            => s_data_in(36,47),
			data_out           => s_data_out(36,47),
			out1               => s_out1(36,47),
			out2               => s_out2(36,47),
			lock_lower_row_out => s_locks_lower_out(36,47),
			lock_lower_row_in  => s_locks_lower_in(36,47),
			in1                => s_in1(36,47),
			in2                => s_in2(36,47),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(47)
		);
	s_in1(36,47)            <= s_out1(37,47);
	s_in2(36,47)            <= s_out2(37,48);
	s_locks_lower_in(36,47) <= s_locks_lower_out(37,47);

		normal_cell_36_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,48),
			fetch              => s_fetch(36,48),
			data_in            => s_data_in(36,48),
			data_out           => s_data_out(36,48),
			out1               => s_out1(36,48),
			out2               => s_out2(36,48),
			lock_lower_row_out => s_locks_lower_out(36,48),
			lock_lower_row_in  => s_locks_lower_in(36,48),
			in1                => s_in1(36,48),
			in2                => s_in2(36,48),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(48)
		);
	s_in1(36,48)            <= s_out1(37,48);
	s_in2(36,48)            <= s_out2(37,49);
	s_locks_lower_in(36,48) <= s_locks_lower_out(37,48);

		normal_cell_36_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,49),
			fetch              => s_fetch(36,49),
			data_in            => s_data_in(36,49),
			data_out           => s_data_out(36,49),
			out1               => s_out1(36,49),
			out2               => s_out2(36,49),
			lock_lower_row_out => s_locks_lower_out(36,49),
			lock_lower_row_in  => s_locks_lower_in(36,49),
			in1                => s_in1(36,49),
			in2                => s_in2(36,49),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(49)
		);
	s_in1(36,49)            <= s_out1(37,49);
	s_in2(36,49)            <= s_out2(37,50);
	s_locks_lower_in(36,49) <= s_locks_lower_out(37,49);

		normal_cell_36_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,50),
			fetch              => s_fetch(36,50),
			data_in            => s_data_in(36,50),
			data_out           => s_data_out(36,50),
			out1               => s_out1(36,50),
			out2               => s_out2(36,50),
			lock_lower_row_out => s_locks_lower_out(36,50),
			lock_lower_row_in  => s_locks_lower_in(36,50),
			in1                => s_in1(36,50),
			in2                => s_in2(36,50),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(50)
		);
	s_in1(36,50)            <= s_out1(37,50);
	s_in2(36,50)            <= s_out2(37,51);
	s_locks_lower_in(36,50) <= s_locks_lower_out(37,50);

		normal_cell_36_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,51),
			fetch              => s_fetch(36,51),
			data_in            => s_data_in(36,51),
			data_out           => s_data_out(36,51),
			out1               => s_out1(36,51),
			out2               => s_out2(36,51),
			lock_lower_row_out => s_locks_lower_out(36,51),
			lock_lower_row_in  => s_locks_lower_in(36,51),
			in1                => s_in1(36,51),
			in2                => s_in2(36,51),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(51)
		);
	s_in1(36,51)            <= s_out1(37,51);
	s_in2(36,51)            <= s_out2(37,52);
	s_locks_lower_in(36,51) <= s_locks_lower_out(37,51);

		normal_cell_36_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,52),
			fetch              => s_fetch(36,52),
			data_in            => s_data_in(36,52),
			data_out           => s_data_out(36,52),
			out1               => s_out1(36,52),
			out2               => s_out2(36,52),
			lock_lower_row_out => s_locks_lower_out(36,52),
			lock_lower_row_in  => s_locks_lower_in(36,52),
			in1                => s_in1(36,52),
			in2                => s_in2(36,52),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(52)
		);
	s_in1(36,52)            <= s_out1(37,52);
	s_in2(36,52)            <= s_out2(37,53);
	s_locks_lower_in(36,52) <= s_locks_lower_out(37,52);

		normal_cell_36_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,53),
			fetch              => s_fetch(36,53),
			data_in            => s_data_in(36,53),
			data_out           => s_data_out(36,53),
			out1               => s_out1(36,53),
			out2               => s_out2(36,53),
			lock_lower_row_out => s_locks_lower_out(36,53),
			lock_lower_row_in  => s_locks_lower_in(36,53),
			in1                => s_in1(36,53),
			in2                => s_in2(36,53),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(53)
		);
	s_in1(36,53)            <= s_out1(37,53);
	s_in2(36,53)            <= s_out2(37,54);
	s_locks_lower_in(36,53) <= s_locks_lower_out(37,53);

		normal_cell_36_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,54),
			fetch              => s_fetch(36,54),
			data_in            => s_data_in(36,54),
			data_out           => s_data_out(36,54),
			out1               => s_out1(36,54),
			out2               => s_out2(36,54),
			lock_lower_row_out => s_locks_lower_out(36,54),
			lock_lower_row_in  => s_locks_lower_in(36,54),
			in1                => s_in1(36,54),
			in2                => s_in2(36,54),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(54)
		);
	s_in1(36,54)            <= s_out1(37,54);
	s_in2(36,54)            <= s_out2(37,55);
	s_locks_lower_in(36,54) <= s_locks_lower_out(37,54);

		normal_cell_36_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,55),
			fetch              => s_fetch(36,55),
			data_in            => s_data_in(36,55),
			data_out           => s_data_out(36,55),
			out1               => s_out1(36,55),
			out2               => s_out2(36,55),
			lock_lower_row_out => s_locks_lower_out(36,55),
			lock_lower_row_in  => s_locks_lower_in(36,55),
			in1                => s_in1(36,55),
			in2                => s_in2(36,55),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(55)
		);
	s_in1(36,55)            <= s_out1(37,55);
	s_in2(36,55)            <= s_out2(37,56);
	s_locks_lower_in(36,55) <= s_locks_lower_out(37,55);

		normal_cell_36_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,56),
			fetch              => s_fetch(36,56),
			data_in            => s_data_in(36,56),
			data_out           => s_data_out(36,56),
			out1               => s_out1(36,56),
			out2               => s_out2(36,56),
			lock_lower_row_out => s_locks_lower_out(36,56),
			lock_lower_row_in  => s_locks_lower_in(36,56),
			in1                => s_in1(36,56),
			in2                => s_in2(36,56),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(56)
		);
	s_in1(36,56)            <= s_out1(37,56);
	s_in2(36,56)            <= s_out2(37,57);
	s_locks_lower_in(36,56) <= s_locks_lower_out(37,56);

		normal_cell_36_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,57),
			fetch              => s_fetch(36,57),
			data_in            => s_data_in(36,57),
			data_out           => s_data_out(36,57),
			out1               => s_out1(36,57),
			out2               => s_out2(36,57),
			lock_lower_row_out => s_locks_lower_out(36,57),
			lock_lower_row_in  => s_locks_lower_in(36,57),
			in1                => s_in1(36,57),
			in2                => s_in2(36,57),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(57)
		);
	s_in1(36,57)            <= s_out1(37,57);
	s_in2(36,57)            <= s_out2(37,58);
	s_locks_lower_in(36,57) <= s_locks_lower_out(37,57);

		normal_cell_36_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,58),
			fetch              => s_fetch(36,58),
			data_in            => s_data_in(36,58),
			data_out           => s_data_out(36,58),
			out1               => s_out1(36,58),
			out2               => s_out2(36,58),
			lock_lower_row_out => s_locks_lower_out(36,58),
			lock_lower_row_in  => s_locks_lower_in(36,58),
			in1                => s_in1(36,58),
			in2                => s_in2(36,58),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(58)
		);
	s_in1(36,58)            <= s_out1(37,58);
	s_in2(36,58)            <= s_out2(37,59);
	s_locks_lower_in(36,58) <= s_locks_lower_out(37,58);

		normal_cell_36_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,59),
			fetch              => s_fetch(36,59),
			data_in            => s_data_in(36,59),
			data_out           => s_data_out(36,59),
			out1               => s_out1(36,59),
			out2               => s_out2(36,59),
			lock_lower_row_out => s_locks_lower_out(36,59),
			lock_lower_row_in  => s_locks_lower_in(36,59),
			in1                => s_in1(36,59),
			in2                => s_in2(36,59),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(59)
		);
	s_in1(36,59)            <= s_out1(37,59);
	s_in2(36,59)            <= s_out2(37,60);
	s_locks_lower_in(36,59) <= s_locks_lower_out(37,59);

		last_col_cell_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(36,60),
			fetch              => s_fetch(36,60),
			data_in            => s_data_in(36,60),
			data_out           => s_data_out(36,60),
			out1               => s_out1(36,60),
			out2               => s_out2(36,60),
			lock_lower_row_out => s_locks_lower_out(36,60),
			lock_lower_row_in  => s_locks_lower_in(36,60),
			in1                => s_in1(36,60),
			in2                => (others => '0'),
			lock_row           => s_locks(36),
			piv_found          => s_piv_found,
			row_data           => s_row_data(36),
			col_data           => s_col_data(60)
		);
	s_in1(36,60)            <= s_out1(37,60);
	s_locks_lower_in(36,60) <= s_locks_lower_out(37,60);

		normal_cell_37_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,1),
			fetch              => s_fetch(37,1),
			data_in            => s_data_in(37,1),
			data_out           => s_data_out(37,1),
			out1               => s_out1(37,1),
			out2               => s_out2(37,1),
			lock_lower_row_out => s_locks_lower_out(37,1),
			lock_lower_row_in  => s_locks_lower_in(37,1),
			in1                => s_in1(37,1),
			in2                => s_in2(37,1),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(1)
		);
	s_in1(37,1)            <= s_out1(38,1);
	s_in2(37,1)            <= s_out2(38,2);
	s_locks_lower_in(37,1) <= s_locks_lower_out(38,1);

		normal_cell_37_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,2),
			fetch              => s_fetch(37,2),
			data_in            => s_data_in(37,2),
			data_out           => s_data_out(37,2),
			out1               => s_out1(37,2),
			out2               => s_out2(37,2),
			lock_lower_row_out => s_locks_lower_out(37,2),
			lock_lower_row_in  => s_locks_lower_in(37,2),
			in1                => s_in1(37,2),
			in2                => s_in2(37,2),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(2)
		);
	s_in1(37,2)            <= s_out1(38,2);
	s_in2(37,2)            <= s_out2(38,3);
	s_locks_lower_in(37,2) <= s_locks_lower_out(38,2);

		normal_cell_37_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,3),
			fetch              => s_fetch(37,3),
			data_in            => s_data_in(37,3),
			data_out           => s_data_out(37,3),
			out1               => s_out1(37,3),
			out2               => s_out2(37,3),
			lock_lower_row_out => s_locks_lower_out(37,3),
			lock_lower_row_in  => s_locks_lower_in(37,3),
			in1                => s_in1(37,3),
			in2                => s_in2(37,3),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(3)
		);
	s_in1(37,3)            <= s_out1(38,3);
	s_in2(37,3)            <= s_out2(38,4);
	s_locks_lower_in(37,3) <= s_locks_lower_out(38,3);

		normal_cell_37_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,4),
			fetch              => s_fetch(37,4),
			data_in            => s_data_in(37,4),
			data_out           => s_data_out(37,4),
			out1               => s_out1(37,4),
			out2               => s_out2(37,4),
			lock_lower_row_out => s_locks_lower_out(37,4),
			lock_lower_row_in  => s_locks_lower_in(37,4),
			in1                => s_in1(37,4),
			in2                => s_in2(37,4),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(4)
		);
	s_in1(37,4)            <= s_out1(38,4);
	s_in2(37,4)            <= s_out2(38,5);
	s_locks_lower_in(37,4) <= s_locks_lower_out(38,4);

		normal_cell_37_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,5),
			fetch              => s_fetch(37,5),
			data_in            => s_data_in(37,5),
			data_out           => s_data_out(37,5),
			out1               => s_out1(37,5),
			out2               => s_out2(37,5),
			lock_lower_row_out => s_locks_lower_out(37,5),
			lock_lower_row_in  => s_locks_lower_in(37,5),
			in1                => s_in1(37,5),
			in2                => s_in2(37,5),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(5)
		);
	s_in1(37,5)            <= s_out1(38,5);
	s_in2(37,5)            <= s_out2(38,6);
	s_locks_lower_in(37,5) <= s_locks_lower_out(38,5);

		normal_cell_37_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,6),
			fetch              => s_fetch(37,6),
			data_in            => s_data_in(37,6),
			data_out           => s_data_out(37,6),
			out1               => s_out1(37,6),
			out2               => s_out2(37,6),
			lock_lower_row_out => s_locks_lower_out(37,6),
			lock_lower_row_in  => s_locks_lower_in(37,6),
			in1                => s_in1(37,6),
			in2                => s_in2(37,6),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(6)
		);
	s_in1(37,6)            <= s_out1(38,6);
	s_in2(37,6)            <= s_out2(38,7);
	s_locks_lower_in(37,6) <= s_locks_lower_out(38,6);

		normal_cell_37_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,7),
			fetch              => s_fetch(37,7),
			data_in            => s_data_in(37,7),
			data_out           => s_data_out(37,7),
			out1               => s_out1(37,7),
			out2               => s_out2(37,7),
			lock_lower_row_out => s_locks_lower_out(37,7),
			lock_lower_row_in  => s_locks_lower_in(37,7),
			in1                => s_in1(37,7),
			in2                => s_in2(37,7),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(7)
		);
	s_in1(37,7)            <= s_out1(38,7);
	s_in2(37,7)            <= s_out2(38,8);
	s_locks_lower_in(37,7) <= s_locks_lower_out(38,7);

		normal_cell_37_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,8),
			fetch              => s_fetch(37,8),
			data_in            => s_data_in(37,8),
			data_out           => s_data_out(37,8),
			out1               => s_out1(37,8),
			out2               => s_out2(37,8),
			lock_lower_row_out => s_locks_lower_out(37,8),
			lock_lower_row_in  => s_locks_lower_in(37,8),
			in1                => s_in1(37,8),
			in2                => s_in2(37,8),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(8)
		);
	s_in1(37,8)            <= s_out1(38,8);
	s_in2(37,8)            <= s_out2(38,9);
	s_locks_lower_in(37,8) <= s_locks_lower_out(38,8);

		normal_cell_37_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,9),
			fetch              => s_fetch(37,9),
			data_in            => s_data_in(37,9),
			data_out           => s_data_out(37,9),
			out1               => s_out1(37,9),
			out2               => s_out2(37,9),
			lock_lower_row_out => s_locks_lower_out(37,9),
			lock_lower_row_in  => s_locks_lower_in(37,9),
			in1                => s_in1(37,9),
			in2                => s_in2(37,9),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(9)
		);
	s_in1(37,9)            <= s_out1(38,9);
	s_in2(37,9)            <= s_out2(38,10);
	s_locks_lower_in(37,9) <= s_locks_lower_out(38,9);

		normal_cell_37_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,10),
			fetch              => s_fetch(37,10),
			data_in            => s_data_in(37,10),
			data_out           => s_data_out(37,10),
			out1               => s_out1(37,10),
			out2               => s_out2(37,10),
			lock_lower_row_out => s_locks_lower_out(37,10),
			lock_lower_row_in  => s_locks_lower_in(37,10),
			in1                => s_in1(37,10),
			in2                => s_in2(37,10),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(10)
		);
	s_in1(37,10)            <= s_out1(38,10);
	s_in2(37,10)            <= s_out2(38,11);
	s_locks_lower_in(37,10) <= s_locks_lower_out(38,10);

		normal_cell_37_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,11),
			fetch              => s_fetch(37,11),
			data_in            => s_data_in(37,11),
			data_out           => s_data_out(37,11),
			out1               => s_out1(37,11),
			out2               => s_out2(37,11),
			lock_lower_row_out => s_locks_lower_out(37,11),
			lock_lower_row_in  => s_locks_lower_in(37,11),
			in1                => s_in1(37,11),
			in2                => s_in2(37,11),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(11)
		);
	s_in1(37,11)            <= s_out1(38,11);
	s_in2(37,11)            <= s_out2(38,12);
	s_locks_lower_in(37,11) <= s_locks_lower_out(38,11);

		normal_cell_37_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,12),
			fetch              => s_fetch(37,12),
			data_in            => s_data_in(37,12),
			data_out           => s_data_out(37,12),
			out1               => s_out1(37,12),
			out2               => s_out2(37,12),
			lock_lower_row_out => s_locks_lower_out(37,12),
			lock_lower_row_in  => s_locks_lower_in(37,12),
			in1                => s_in1(37,12),
			in2                => s_in2(37,12),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(12)
		);
	s_in1(37,12)            <= s_out1(38,12);
	s_in2(37,12)            <= s_out2(38,13);
	s_locks_lower_in(37,12) <= s_locks_lower_out(38,12);

		normal_cell_37_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,13),
			fetch              => s_fetch(37,13),
			data_in            => s_data_in(37,13),
			data_out           => s_data_out(37,13),
			out1               => s_out1(37,13),
			out2               => s_out2(37,13),
			lock_lower_row_out => s_locks_lower_out(37,13),
			lock_lower_row_in  => s_locks_lower_in(37,13),
			in1                => s_in1(37,13),
			in2                => s_in2(37,13),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(13)
		);
	s_in1(37,13)            <= s_out1(38,13);
	s_in2(37,13)            <= s_out2(38,14);
	s_locks_lower_in(37,13) <= s_locks_lower_out(38,13);

		normal_cell_37_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,14),
			fetch              => s_fetch(37,14),
			data_in            => s_data_in(37,14),
			data_out           => s_data_out(37,14),
			out1               => s_out1(37,14),
			out2               => s_out2(37,14),
			lock_lower_row_out => s_locks_lower_out(37,14),
			lock_lower_row_in  => s_locks_lower_in(37,14),
			in1                => s_in1(37,14),
			in2                => s_in2(37,14),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(14)
		);
	s_in1(37,14)            <= s_out1(38,14);
	s_in2(37,14)            <= s_out2(38,15);
	s_locks_lower_in(37,14) <= s_locks_lower_out(38,14);

		normal_cell_37_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,15),
			fetch              => s_fetch(37,15),
			data_in            => s_data_in(37,15),
			data_out           => s_data_out(37,15),
			out1               => s_out1(37,15),
			out2               => s_out2(37,15),
			lock_lower_row_out => s_locks_lower_out(37,15),
			lock_lower_row_in  => s_locks_lower_in(37,15),
			in1                => s_in1(37,15),
			in2                => s_in2(37,15),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(15)
		);
	s_in1(37,15)            <= s_out1(38,15);
	s_in2(37,15)            <= s_out2(38,16);
	s_locks_lower_in(37,15) <= s_locks_lower_out(38,15);

		normal_cell_37_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,16),
			fetch              => s_fetch(37,16),
			data_in            => s_data_in(37,16),
			data_out           => s_data_out(37,16),
			out1               => s_out1(37,16),
			out2               => s_out2(37,16),
			lock_lower_row_out => s_locks_lower_out(37,16),
			lock_lower_row_in  => s_locks_lower_in(37,16),
			in1                => s_in1(37,16),
			in2                => s_in2(37,16),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(16)
		);
	s_in1(37,16)            <= s_out1(38,16);
	s_in2(37,16)            <= s_out2(38,17);
	s_locks_lower_in(37,16) <= s_locks_lower_out(38,16);

		normal_cell_37_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,17),
			fetch              => s_fetch(37,17),
			data_in            => s_data_in(37,17),
			data_out           => s_data_out(37,17),
			out1               => s_out1(37,17),
			out2               => s_out2(37,17),
			lock_lower_row_out => s_locks_lower_out(37,17),
			lock_lower_row_in  => s_locks_lower_in(37,17),
			in1                => s_in1(37,17),
			in2                => s_in2(37,17),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(17)
		);
	s_in1(37,17)            <= s_out1(38,17);
	s_in2(37,17)            <= s_out2(38,18);
	s_locks_lower_in(37,17) <= s_locks_lower_out(38,17);

		normal_cell_37_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,18),
			fetch              => s_fetch(37,18),
			data_in            => s_data_in(37,18),
			data_out           => s_data_out(37,18),
			out1               => s_out1(37,18),
			out2               => s_out2(37,18),
			lock_lower_row_out => s_locks_lower_out(37,18),
			lock_lower_row_in  => s_locks_lower_in(37,18),
			in1                => s_in1(37,18),
			in2                => s_in2(37,18),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(18)
		);
	s_in1(37,18)            <= s_out1(38,18);
	s_in2(37,18)            <= s_out2(38,19);
	s_locks_lower_in(37,18) <= s_locks_lower_out(38,18);

		normal_cell_37_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,19),
			fetch              => s_fetch(37,19),
			data_in            => s_data_in(37,19),
			data_out           => s_data_out(37,19),
			out1               => s_out1(37,19),
			out2               => s_out2(37,19),
			lock_lower_row_out => s_locks_lower_out(37,19),
			lock_lower_row_in  => s_locks_lower_in(37,19),
			in1                => s_in1(37,19),
			in2                => s_in2(37,19),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(19)
		);
	s_in1(37,19)            <= s_out1(38,19);
	s_in2(37,19)            <= s_out2(38,20);
	s_locks_lower_in(37,19) <= s_locks_lower_out(38,19);

		normal_cell_37_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,20),
			fetch              => s_fetch(37,20),
			data_in            => s_data_in(37,20),
			data_out           => s_data_out(37,20),
			out1               => s_out1(37,20),
			out2               => s_out2(37,20),
			lock_lower_row_out => s_locks_lower_out(37,20),
			lock_lower_row_in  => s_locks_lower_in(37,20),
			in1                => s_in1(37,20),
			in2                => s_in2(37,20),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(20)
		);
	s_in1(37,20)            <= s_out1(38,20);
	s_in2(37,20)            <= s_out2(38,21);
	s_locks_lower_in(37,20) <= s_locks_lower_out(38,20);

		normal_cell_37_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,21),
			fetch              => s_fetch(37,21),
			data_in            => s_data_in(37,21),
			data_out           => s_data_out(37,21),
			out1               => s_out1(37,21),
			out2               => s_out2(37,21),
			lock_lower_row_out => s_locks_lower_out(37,21),
			lock_lower_row_in  => s_locks_lower_in(37,21),
			in1                => s_in1(37,21),
			in2                => s_in2(37,21),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(21)
		);
	s_in1(37,21)            <= s_out1(38,21);
	s_in2(37,21)            <= s_out2(38,22);
	s_locks_lower_in(37,21) <= s_locks_lower_out(38,21);

		normal_cell_37_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,22),
			fetch              => s_fetch(37,22),
			data_in            => s_data_in(37,22),
			data_out           => s_data_out(37,22),
			out1               => s_out1(37,22),
			out2               => s_out2(37,22),
			lock_lower_row_out => s_locks_lower_out(37,22),
			lock_lower_row_in  => s_locks_lower_in(37,22),
			in1                => s_in1(37,22),
			in2                => s_in2(37,22),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(22)
		);
	s_in1(37,22)            <= s_out1(38,22);
	s_in2(37,22)            <= s_out2(38,23);
	s_locks_lower_in(37,22) <= s_locks_lower_out(38,22);

		normal_cell_37_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,23),
			fetch              => s_fetch(37,23),
			data_in            => s_data_in(37,23),
			data_out           => s_data_out(37,23),
			out1               => s_out1(37,23),
			out2               => s_out2(37,23),
			lock_lower_row_out => s_locks_lower_out(37,23),
			lock_lower_row_in  => s_locks_lower_in(37,23),
			in1                => s_in1(37,23),
			in2                => s_in2(37,23),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(23)
		);
	s_in1(37,23)            <= s_out1(38,23);
	s_in2(37,23)            <= s_out2(38,24);
	s_locks_lower_in(37,23) <= s_locks_lower_out(38,23);

		normal_cell_37_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,24),
			fetch              => s_fetch(37,24),
			data_in            => s_data_in(37,24),
			data_out           => s_data_out(37,24),
			out1               => s_out1(37,24),
			out2               => s_out2(37,24),
			lock_lower_row_out => s_locks_lower_out(37,24),
			lock_lower_row_in  => s_locks_lower_in(37,24),
			in1                => s_in1(37,24),
			in2                => s_in2(37,24),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(24)
		);
	s_in1(37,24)            <= s_out1(38,24);
	s_in2(37,24)            <= s_out2(38,25);
	s_locks_lower_in(37,24) <= s_locks_lower_out(38,24);

		normal_cell_37_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,25),
			fetch              => s_fetch(37,25),
			data_in            => s_data_in(37,25),
			data_out           => s_data_out(37,25),
			out1               => s_out1(37,25),
			out2               => s_out2(37,25),
			lock_lower_row_out => s_locks_lower_out(37,25),
			lock_lower_row_in  => s_locks_lower_in(37,25),
			in1                => s_in1(37,25),
			in2                => s_in2(37,25),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(25)
		);
	s_in1(37,25)            <= s_out1(38,25);
	s_in2(37,25)            <= s_out2(38,26);
	s_locks_lower_in(37,25) <= s_locks_lower_out(38,25);

		normal_cell_37_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,26),
			fetch              => s_fetch(37,26),
			data_in            => s_data_in(37,26),
			data_out           => s_data_out(37,26),
			out1               => s_out1(37,26),
			out2               => s_out2(37,26),
			lock_lower_row_out => s_locks_lower_out(37,26),
			lock_lower_row_in  => s_locks_lower_in(37,26),
			in1                => s_in1(37,26),
			in2                => s_in2(37,26),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(26)
		);
	s_in1(37,26)            <= s_out1(38,26);
	s_in2(37,26)            <= s_out2(38,27);
	s_locks_lower_in(37,26) <= s_locks_lower_out(38,26);

		normal_cell_37_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,27),
			fetch              => s_fetch(37,27),
			data_in            => s_data_in(37,27),
			data_out           => s_data_out(37,27),
			out1               => s_out1(37,27),
			out2               => s_out2(37,27),
			lock_lower_row_out => s_locks_lower_out(37,27),
			lock_lower_row_in  => s_locks_lower_in(37,27),
			in1                => s_in1(37,27),
			in2                => s_in2(37,27),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(27)
		);
	s_in1(37,27)            <= s_out1(38,27);
	s_in2(37,27)            <= s_out2(38,28);
	s_locks_lower_in(37,27) <= s_locks_lower_out(38,27);

		normal_cell_37_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,28),
			fetch              => s_fetch(37,28),
			data_in            => s_data_in(37,28),
			data_out           => s_data_out(37,28),
			out1               => s_out1(37,28),
			out2               => s_out2(37,28),
			lock_lower_row_out => s_locks_lower_out(37,28),
			lock_lower_row_in  => s_locks_lower_in(37,28),
			in1                => s_in1(37,28),
			in2                => s_in2(37,28),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(28)
		);
	s_in1(37,28)            <= s_out1(38,28);
	s_in2(37,28)            <= s_out2(38,29);
	s_locks_lower_in(37,28) <= s_locks_lower_out(38,28);

		normal_cell_37_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,29),
			fetch              => s_fetch(37,29),
			data_in            => s_data_in(37,29),
			data_out           => s_data_out(37,29),
			out1               => s_out1(37,29),
			out2               => s_out2(37,29),
			lock_lower_row_out => s_locks_lower_out(37,29),
			lock_lower_row_in  => s_locks_lower_in(37,29),
			in1                => s_in1(37,29),
			in2                => s_in2(37,29),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(29)
		);
	s_in1(37,29)            <= s_out1(38,29);
	s_in2(37,29)            <= s_out2(38,30);
	s_locks_lower_in(37,29) <= s_locks_lower_out(38,29);

		normal_cell_37_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,30),
			fetch              => s_fetch(37,30),
			data_in            => s_data_in(37,30),
			data_out           => s_data_out(37,30),
			out1               => s_out1(37,30),
			out2               => s_out2(37,30),
			lock_lower_row_out => s_locks_lower_out(37,30),
			lock_lower_row_in  => s_locks_lower_in(37,30),
			in1                => s_in1(37,30),
			in2                => s_in2(37,30),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(30)
		);
	s_in1(37,30)            <= s_out1(38,30);
	s_in2(37,30)            <= s_out2(38,31);
	s_locks_lower_in(37,30) <= s_locks_lower_out(38,30);

		normal_cell_37_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,31),
			fetch              => s_fetch(37,31),
			data_in            => s_data_in(37,31),
			data_out           => s_data_out(37,31),
			out1               => s_out1(37,31),
			out2               => s_out2(37,31),
			lock_lower_row_out => s_locks_lower_out(37,31),
			lock_lower_row_in  => s_locks_lower_in(37,31),
			in1                => s_in1(37,31),
			in2                => s_in2(37,31),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(31)
		);
	s_in1(37,31)            <= s_out1(38,31);
	s_in2(37,31)            <= s_out2(38,32);
	s_locks_lower_in(37,31) <= s_locks_lower_out(38,31);

		normal_cell_37_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,32),
			fetch              => s_fetch(37,32),
			data_in            => s_data_in(37,32),
			data_out           => s_data_out(37,32),
			out1               => s_out1(37,32),
			out2               => s_out2(37,32),
			lock_lower_row_out => s_locks_lower_out(37,32),
			lock_lower_row_in  => s_locks_lower_in(37,32),
			in1                => s_in1(37,32),
			in2                => s_in2(37,32),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(32)
		);
	s_in1(37,32)            <= s_out1(38,32);
	s_in2(37,32)            <= s_out2(38,33);
	s_locks_lower_in(37,32) <= s_locks_lower_out(38,32);

		normal_cell_37_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,33),
			fetch              => s_fetch(37,33),
			data_in            => s_data_in(37,33),
			data_out           => s_data_out(37,33),
			out1               => s_out1(37,33),
			out2               => s_out2(37,33),
			lock_lower_row_out => s_locks_lower_out(37,33),
			lock_lower_row_in  => s_locks_lower_in(37,33),
			in1                => s_in1(37,33),
			in2                => s_in2(37,33),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(33)
		);
	s_in1(37,33)            <= s_out1(38,33);
	s_in2(37,33)            <= s_out2(38,34);
	s_locks_lower_in(37,33) <= s_locks_lower_out(38,33);

		normal_cell_37_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,34),
			fetch              => s_fetch(37,34),
			data_in            => s_data_in(37,34),
			data_out           => s_data_out(37,34),
			out1               => s_out1(37,34),
			out2               => s_out2(37,34),
			lock_lower_row_out => s_locks_lower_out(37,34),
			lock_lower_row_in  => s_locks_lower_in(37,34),
			in1                => s_in1(37,34),
			in2                => s_in2(37,34),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(34)
		);
	s_in1(37,34)            <= s_out1(38,34);
	s_in2(37,34)            <= s_out2(38,35);
	s_locks_lower_in(37,34) <= s_locks_lower_out(38,34);

		normal_cell_37_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,35),
			fetch              => s_fetch(37,35),
			data_in            => s_data_in(37,35),
			data_out           => s_data_out(37,35),
			out1               => s_out1(37,35),
			out2               => s_out2(37,35),
			lock_lower_row_out => s_locks_lower_out(37,35),
			lock_lower_row_in  => s_locks_lower_in(37,35),
			in1                => s_in1(37,35),
			in2                => s_in2(37,35),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(35)
		);
	s_in1(37,35)            <= s_out1(38,35);
	s_in2(37,35)            <= s_out2(38,36);
	s_locks_lower_in(37,35) <= s_locks_lower_out(38,35);

		normal_cell_37_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,36),
			fetch              => s_fetch(37,36),
			data_in            => s_data_in(37,36),
			data_out           => s_data_out(37,36),
			out1               => s_out1(37,36),
			out2               => s_out2(37,36),
			lock_lower_row_out => s_locks_lower_out(37,36),
			lock_lower_row_in  => s_locks_lower_in(37,36),
			in1                => s_in1(37,36),
			in2                => s_in2(37,36),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(36)
		);
	s_in1(37,36)            <= s_out1(38,36);
	s_in2(37,36)            <= s_out2(38,37);
	s_locks_lower_in(37,36) <= s_locks_lower_out(38,36);

		normal_cell_37_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,37),
			fetch              => s_fetch(37,37),
			data_in            => s_data_in(37,37),
			data_out           => s_data_out(37,37),
			out1               => s_out1(37,37),
			out2               => s_out2(37,37),
			lock_lower_row_out => s_locks_lower_out(37,37),
			lock_lower_row_in  => s_locks_lower_in(37,37),
			in1                => s_in1(37,37),
			in2                => s_in2(37,37),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(37)
		);
	s_in1(37,37)            <= s_out1(38,37);
	s_in2(37,37)            <= s_out2(38,38);
	s_locks_lower_in(37,37) <= s_locks_lower_out(38,37);

		normal_cell_37_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,38),
			fetch              => s_fetch(37,38),
			data_in            => s_data_in(37,38),
			data_out           => s_data_out(37,38),
			out1               => s_out1(37,38),
			out2               => s_out2(37,38),
			lock_lower_row_out => s_locks_lower_out(37,38),
			lock_lower_row_in  => s_locks_lower_in(37,38),
			in1                => s_in1(37,38),
			in2                => s_in2(37,38),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(38)
		);
	s_in1(37,38)            <= s_out1(38,38);
	s_in2(37,38)            <= s_out2(38,39);
	s_locks_lower_in(37,38) <= s_locks_lower_out(38,38);

		normal_cell_37_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,39),
			fetch              => s_fetch(37,39),
			data_in            => s_data_in(37,39),
			data_out           => s_data_out(37,39),
			out1               => s_out1(37,39),
			out2               => s_out2(37,39),
			lock_lower_row_out => s_locks_lower_out(37,39),
			lock_lower_row_in  => s_locks_lower_in(37,39),
			in1                => s_in1(37,39),
			in2                => s_in2(37,39),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(39)
		);
	s_in1(37,39)            <= s_out1(38,39);
	s_in2(37,39)            <= s_out2(38,40);
	s_locks_lower_in(37,39) <= s_locks_lower_out(38,39);

		normal_cell_37_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,40),
			fetch              => s_fetch(37,40),
			data_in            => s_data_in(37,40),
			data_out           => s_data_out(37,40),
			out1               => s_out1(37,40),
			out2               => s_out2(37,40),
			lock_lower_row_out => s_locks_lower_out(37,40),
			lock_lower_row_in  => s_locks_lower_in(37,40),
			in1                => s_in1(37,40),
			in2                => s_in2(37,40),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(40)
		);
	s_in1(37,40)            <= s_out1(38,40);
	s_in2(37,40)            <= s_out2(38,41);
	s_locks_lower_in(37,40) <= s_locks_lower_out(38,40);

		normal_cell_37_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,41),
			fetch              => s_fetch(37,41),
			data_in            => s_data_in(37,41),
			data_out           => s_data_out(37,41),
			out1               => s_out1(37,41),
			out2               => s_out2(37,41),
			lock_lower_row_out => s_locks_lower_out(37,41),
			lock_lower_row_in  => s_locks_lower_in(37,41),
			in1                => s_in1(37,41),
			in2                => s_in2(37,41),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(41)
		);
	s_in1(37,41)            <= s_out1(38,41);
	s_in2(37,41)            <= s_out2(38,42);
	s_locks_lower_in(37,41) <= s_locks_lower_out(38,41);

		normal_cell_37_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,42),
			fetch              => s_fetch(37,42),
			data_in            => s_data_in(37,42),
			data_out           => s_data_out(37,42),
			out1               => s_out1(37,42),
			out2               => s_out2(37,42),
			lock_lower_row_out => s_locks_lower_out(37,42),
			lock_lower_row_in  => s_locks_lower_in(37,42),
			in1                => s_in1(37,42),
			in2                => s_in2(37,42),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(42)
		);
	s_in1(37,42)            <= s_out1(38,42);
	s_in2(37,42)            <= s_out2(38,43);
	s_locks_lower_in(37,42) <= s_locks_lower_out(38,42);

		normal_cell_37_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,43),
			fetch              => s_fetch(37,43),
			data_in            => s_data_in(37,43),
			data_out           => s_data_out(37,43),
			out1               => s_out1(37,43),
			out2               => s_out2(37,43),
			lock_lower_row_out => s_locks_lower_out(37,43),
			lock_lower_row_in  => s_locks_lower_in(37,43),
			in1                => s_in1(37,43),
			in2                => s_in2(37,43),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(43)
		);
	s_in1(37,43)            <= s_out1(38,43);
	s_in2(37,43)            <= s_out2(38,44);
	s_locks_lower_in(37,43) <= s_locks_lower_out(38,43);

		normal_cell_37_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,44),
			fetch              => s_fetch(37,44),
			data_in            => s_data_in(37,44),
			data_out           => s_data_out(37,44),
			out1               => s_out1(37,44),
			out2               => s_out2(37,44),
			lock_lower_row_out => s_locks_lower_out(37,44),
			lock_lower_row_in  => s_locks_lower_in(37,44),
			in1                => s_in1(37,44),
			in2                => s_in2(37,44),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(44)
		);
	s_in1(37,44)            <= s_out1(38,44);
	s_in2(37,44)            <= s_out2(38,45);
	s_locks_lower_in(37,44) <= s_locks_lower_out(38,44);

		normal_cell_37_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,45),
			fetch              => s_fetch(37,45),
			data_in            => s_data_in(37,45),
			data_out           => s_data_out(37,45),
			out1               => s_out1(37,45),
			out2               => s_out2(37,45),
			lock_lower_row_out => s_locks_lower_out(37,45),
			lock_lower_row_in  => s_locks_lower_in(37,45),
			in1                => s_in1(37,45),
			in2                => s_in2(37,45),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(45)
		);
	s_in1(37,45)            <= s_out1(38,45);
	s_in2(37,45)            <= s_out2(38,46);
	s_locks_lower_in(37,45) <= s_locks_lower_out(38,45);

		normal_cell_37_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,46),
			fetch              => s_fetch(37,46),
			data_in            => s_data_in(37,46),
			data_out           => s_data_out(37,46),
			out1               => s_out1(37,46),
			out2               => s_out2(37,46),
			lock_lower_row_out => s_locks_lower_out(37,46),
			lock_lower_row_in  => s_locks_lower_in(37,46),
			in1                => s_in1(37,46),
			in2                => s_in2(37,46),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(46)
		);
	s_in1(37,46)            <= s_out1(38,46);
	s_in2(37,46)            <= s_out2(38,47);
	s_locks_lower_in(37,46) <= s_locks_lower_out(38,46);

		normal_cell_37_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,47),
			fetch              => s_fetch(37,47),
			data_in            => s_data_in(37,47),
			data_out           => s_data_out(37,47),
			out1               => s_out1(37,47),
			out2               => s_out2(37,47),
			lock_lower_row_out => s_locks_lower_out(37,47),
			lock_lower_row_in  => s_locks_lower_in(37,47),
			in1                => s_in1(37,47),
			in2                => s_in2(37,47),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(47)
		);
	s_in1(37,47)            <= s_out1(38,47);
	s_in2(37,47)            <= s_out2(38,48);
	s_locks_lower_in(37,47) <= s_locks_lower_out(38,47);

		normal_cell_37_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,48),
			fetch              => s_fetch(37,48),
			data_in            => s_data_in(37,48),
			data_out           => s_data_out(37,48),
			out1               => s_out1(37,48),
			out2               => s_out2(37,48),
			lock_lower_row_out => s_locks_lower_out(37,48),
			lock_lower_row_in  => s_locks_lower_in(37,48),
			in1                => s_in1(37,48),
			in2                => s_in2(37,48),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(48)
		);
	s_in1(37,48)            <= s_out1(38,48);
	s_in2(37,48)            <= s_out2(38,49);
	s_locks_lower_in(37,48) <= s_locks_lower_out(38,48);

		normal_cell_37_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,49),
			fetch              => s_fetch(37,49),
			data_in            => s_data_in(37,49),
			data_out           => s_data_out(37,49),
			out1               => s_out1(37,49),
			out2               => s_out2(37,49),
			lock_lower_row_out => s_locks_lower_out(37,49),
			lock_lower_row_in  => s_locks_lower_in(37,49),
			in1                => s_in1(37,49),
			in2                => s_in2(37,49),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(49)
		);
	s_in1(37,49)            <= s_out1(38,49);
	s_in2(37,49)            <= s_out2(38,50);
	s_locks_lower_in(37,49) <= s_locks_lower_out(38,49);

		normal_cell_37_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,50),
			fetch              => s_fetch(37,50),
			data_in            => s_data_in(37,50),
			data_out           => s_data_out(37,50),
			out1               => s_out1(37,50),
			out2               => s_out2(37,50),
			lock_lower_row_out => s_locks_lower_out(37,50),
			lock_lower_row_in  => s_locks_lower_in(37,50),
			in1                => s_in1(37,50),
			in2                => s_in2(37,50),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(50)
		);
	s_in1(37,50)            <= s_out1(38,50);
	s_in2(37,50)            <= s_out2(38,51);
	s_locks_lower_in(37,50) <= s_locks_lower_out(38,50);

		normal_cell_37_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,51),
			fetch              => s_fetch(37,51),
			data_in            => s_data_in(37,51),
			data_out           => s_data_out(37,51),
			out1               => s_out1(37,51),
			out2               => s_out2(37,51),
			lock_lower_row_out => s_locks_lower_out(37,51),
			lock_lower_row_in  => s_locks_lower_in(37,51),
			in1                => s_in1(37,51),
			in2                => s_in2(37,51),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(51)
		);
	s_in1(37,51)            <= s_out1(38,51);
	s_in2(37,51)            <= s_out2(38,52);
	s_locks_lower_in(37,51) <= s_locks_lower_out(38,51);

		normal_cell_37_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,52),
			fetch              => s_fetch(37,52),
			data_in            => s_data_in(37,52),
			data_out           => s_data_out(37,52),
			out1               => s_out1(37,52),
			out2               => s_out2(37,52),
			lock_lower_row_out => s_locks_lower_out(37,52),
			lock_lower_row_in  => s_locks_lower_in(37,52),
			in1                => s_in1(37,52),
			in2                => s_in2(37,52),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(52)
		);
	s_in1(37,52)            <= s_out1(38,52);
	s_in2(37,52)            <= s_out2(38,53);
	s_locks_lower_in(37,52) <= s_locks_lower_out(38,52);

		normal_cell_37_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,53),
			fetch              => s_fetch(37,53),
			data_in            => s_data_in(37,53),
			data_out           => s_data_out(37,53),
			out1               => s_out1(37,53),
			out2               => s_out2(37,53),
			lock_lower_row_out => s_locks_lower_out(37,53),
			lock_lower_row_in  => s_locks_lower_in(37,53),
			in1                => s_in1(37,53),
			in2                => s_in2(37,53),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(53)
		);
	s_in1(37,53)            <= s_out1(38,53);
	s_in2(37,53)            <= s_out2(38,54);
	s_locks_lower_in(37,53) <= s_locks_lower_out(38,53);

		normal_cell_37_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,54),
			fetch              => s_fetch(37,54),
			data_in            => s_data_in(37,54),
			data_out           => s_data_out(37,54),
			out1               => s_out1(37,54),
			out2               => s_out2(37,54),
			lock_lower_row_out => s_locks_lower_out(37,54),
			lock_lower_row_in  => s_locks_lower_in(37,54),
			in1                => s_in1(37,54),
			in2                => s_in2(37,54),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(54)
		);
	s_in1(37,54)            <= s_out1(38,54);
	s_in2(37,54)            <= s_out2(38,55);
	s_locks_lower_in(37,54) <= s_locks_lower_out(38,54);

		normal_cell_37_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,55),
			fetch              => s_fetch(37,55),
			data_in            => s_data_in(37,55),
			data_out           => s_data_out(37,55),
			out1               => s_out1(37,55),
			out2               => s_out2(37,55),
			lock_lower_row_out => s_locks_lower_out(37,55),
			lock_lower_row_in  => s_locks_lower_in(37,55),
			in1                => s_in1(37,55),
			in2                => s_in2(37,55),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(55)
		);
	s_in1(37,55)            <= s_out1(38,55);
	s_in2(37,55)            <= s_out2(38,56);
	s_locks_lower_in(37,55) <= s_locks_lower_out(38,55);

		normal_cell_37_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,56),
			fetch              => s_fetch(37,56),
			data_in            => s_data_in(37,56),
			data_out           => s_data_out(37,56),
			out1               => s_out1(37,56),
			out2               => s_out2(37,56),
			lock_lower_row_out => s_locks_lower_out(37,56),
			lock_lower_row_in  => s_locks_lower_in(37,56),
			in1                => s_in1(37,56),
			in2                => s_in2(37,56),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(56)
		);
	s_in1(37,56)            <= s_out1(38,56);
	s_in2(37,56)            <= s_out2(38,57);
	s_locks_lower_in(37,56) <= s_locks_lower_out(38,56);

		normal_cell_37_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,57),
			fetch              => s_fetch(37,57),
			data_in            => s_data_in(37,57),
			data_out           => s_data_out(37,57),
			out1               => s_out1(37,57),
			out2               => s_out2(37,57),
			lock_lower_row_out => s_locks_lower_out(37,57),
			lock_lower_row_in  => s_locks_lower_in(37,57),
			in1                => s_in1(37,57),
			in2                => s_in2(37,57),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(57)
		);
	s_in1(37,57)            <= s_out1(38,57);
	s_in2(37,57)            <= s_out2(38,58);
	s_locks_lower_in(37,57) <= s_locks_lower_out(38,57);

		normal_cell_37_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,58),
			fetch              => s_fetch(37,58),
			data_in            => s_data_in(37,58),
			data_out           => s_data_out(37,58),
			out1               => s_out1(37,58),
			out2               => s_out2(37,58),
			lock_lower_row_out => s_locks_lower_out(37,58),
			lock_lower_row_in  => s_locks_lower_in(37,58),
			in1                => s_in1(37,58),
			in2                => s_in2(37,58),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(58)
		);
	s_in1(37,58)            <= s_out1(38,58);
	s_in2(37,58)            <= s_out2(38,59);
	s_locks_lower_in(37,58) <= s_locks_lower_out(38,58);

		normal_cell_37_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,59),
			fetch              => s_fetch(37,59),
			data_in            => s_data_in(37,59),
			data_out           => s_data_out(37,59),
			out1               => s_out1(37,59),
			out2               => s_out2(37,59),
			lock_lower_row_out => s_locks_lower_out(37,59),
			lock_lower_row_in  => s_locks_lower_in(37,59),
			in1                => s_in1(37,59),
			in2                => s_in2(37,59),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(59)
		);
	s_in1(37,59)            <= s_out1(38,59);
	s_in2(37,59)            <= s_out2(38,60);
	s_locks_lower_in(37,59) <= s_locks_lower_out(38,59);

		last_col_cell_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(37,60),
			fetch              => s_fetch(37,60),
			data_in            => s_data_in(37,60),
			data_out           => s_data_out(37,60),
			out1               => s_out1(37,60),
			out2               => s_out2(37,60),
			lock_lower_row_out => s_locks_lower_out(37,60),
			lock_lower_row_in  => s_locks_lower_in(37,60),
			in1                => s_in1(37,60),
			in2                => (others => '0'),
			lock_row           => s_locks(37),
			piv_found          => s_piv_found,
			row_data           => s_row_data(37),
			col_data           => s_col_data(60)
		);
	s_in1(37,60)            <= s_out1(38,60);
	s_locks_lower_in(37,60) <= s_locks_lower_out(38,60);

		normal_cell_38_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,1),
			fetch              => s_fetch(38,1),
			data_in            => s_data_in(38,1),
			data_out           => s_data_out(38,1),
			out1               => s_out1(38,1),
			out2               => s_out2(38,1),
			lock_lower_row_out => s_locks_lower_out(38,1),
			lock_lower_row_in  => s_locks_lower_in(38,1),
			in1                => s_in1(38,1),
			in2                => s_in2(38,1),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(1)
		);
	s_in1(38,1)            <= s_out1(39,1);
	s_in2(38,1)            <= s_out2(39,2);
	s_locks_lower_in(38,1) <= s_locks_lower_out(39,1);

		normal_cell_38_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,2),
			fetch              => s_fetch(38,2),
			data_in            => s_data_in(38,2),
			data_out           => s_data_out(38,2),
			out1               => s_out1(38,2),
			out2               => s_out2(38,2),
			lock_lower_row_out => s_locks_lower_out(38,2),
			lock_lower_row_in  => s_locks_lower_in(38,2),
			in1                => s_in1(38,2),
			in2                => s_in2(38,2),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(2)
		);
	s_in1(38,2)            <= s_out1(39,2);
	s_in2(38,2)            <= s_out2(39,3);
	s_locks_lower_in(38,2) <= s_locks_lower_out(39,2);

		normal_cell_38_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,3),
			fetch              => s_fetch(38,3),
			data_in            => s_data_in(38,3),
			data_out           => s_data_out(38,3),
			out1               => s_out1(38,3),
			out2               => s_out2(38,3),
			lock_lower_row_out => s_locks_lower_out(38,3),
			lock_lower_row_in  => s_locks_lower_in(38,3),
			in1                => s_in1(38,3),
			in2                => s_in2(38,3),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(3)
		);
	s_in1(38,3)            <= s_out1(39,3);
	s_in2(38,3)            <= s_out2(39,4);
	s_locks_lower_in(38,3) <= s_locks_lower_out(39,3);

		normal_cell_38_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,4),
			fetch              => s_fetch(38,4),
			data_in            => s_data_in(38,4),
			data_out           => s_data_out(38,4),
			out1               => s_out1(38,4),
			out2               => s_out2(38,4),
			lock_lower_row_out => s_locks_lower_out(38,4),
			lock_lower_row_in  => s_locks_lower_in(38,4),
			in1                => s_in1(38,4),
			in2                => s_in2(38,4),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(4)
		);
	s_in1(38,4)            <= s_out1(39,4);
	s_in2(38,4)            <= s_out2(39,5);
	s_locks_lower_in(38,4) <= s_locks_lower_out(39,4);

		normal_cell_38_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,5),
			fetch              => s_fetch(38,5),
			data_in            => s_data_in(38,5),
			data_out           => s_data_out(38,5),
			out1               => s_out1(38,5),
			out2               => s_out2(38,5),
			lock_lower_row_out => s_locks_lower_out(38,5),
			lock_lower_row_in  => s_locks_lower_in(38,5),
			in1                => s_in1(38,5),
			in2                => s_in2(38,5),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(5)
		);
	s_in1(38,5)            <= s_out1(39,5);
	s_in2(38,5)            <= s_out2(39,6);
	s_locks_lower_in(38,5) <= s_locks_lower_out(39,5);

		normal_cell_38_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,6),
			fetch              => s_fetch(38,6),
			data_in            => s_data_in(38,6),
			data_out           => s_data_out(38,6),
			out1               => s_out1(38,6),
			out2               => s_out2(38,6),
			lock_lower_row_out => s_locks_lower_out(38,6),
			lock_lower_row_in  => s_locks_lower_in(38,6),
			in1                => s_in1(38,6),
			in2                => s_in2(38,6),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(6)
		);
	s_in1(38,6)            <= s_out1(39,6);
	s_in2(38,6)            <= s_out2(39,7);
	s_locks_lower_in(38,6) <= s_locks_lower_out(39,6);

		normal_cell_38_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,7),
			fetch              => s_fetch(38,7),
			data_in            => s_data_in(38,7),
			data_out           => s_data_out(38,7),
			out1               => s_out1(38,7),
			out2               => s_out2(38,7),
			lock_lower_row_out => s_locks_lower_out(38,7),
			lock_lower_row_in  => s_locks_lower_in(38,7),
			in1                => s_in1(38,7),
			in2                => s_in2(38,7),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(7)
		);
	s_in1(38,7)            <= s_out1(39,7);
	s_in2(38,7)            <= s_out2(39,8);
	s_locks_lower_in(38,7) <= s_locks_lower_out(39,7);

		normal_cell_38_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,8),
			fetch              => s_fetch(38,8),
			data_in            => s_data_in(38,8),
			data_out           => s_data_out(38,8),
			out1               => s_out1(38,8),
			out2               => s_out2(38,8),
			lock_lower_row_out => s_locks_lower_out(38,8),
			lock_lower_row_in  => s_locks_lower_in(38,8),
			in1                => s_in1(38,8),
			in2                => s_in2(38,8),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(8)
		);
	s_in1(38,8)            <= s_out1(39,8);
	s_in2(38,8)            <= s_out2(39,9);
	s_locks_lower_in(38,8) <= s_locks_lower_out(39,8);

		normal_cell_38_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,9),
			fetch              => s_fetch(38,9),
			data_in            => s_data_in(38,9),
			data_out           => s_data_out(38,9),
			out1               => s_out1(38,9),
			out2               => s_out2(38,9),
			lock_lower_row_out => s_locks_lower_out(38,9),
			lock_lower_row_in  => s_locks_lower_in(38,9),
			in1                => s_in1(38,9),
			in2                => s_in2(38,9),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(9)
		);
	s_in1(38,9)            <= s_out1(39,9);
	s_in2(38,9)            <= s_out2(39,10);
	s_locks_lower_in(38,9) <= s_locks_lower_out(39,9);

		normal_cell_38_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,10),
			fetch              => s_fetch(38,10),
			data_in            => s_data_in(38,10),
			data_out           => s_data_out(38,10),
			out1               => s_out1(38,10),
			out2               => s_out2(38,10),
			lock_lower_row_out => s_locks_lower_out(38,10),
			lock_lower_row_in  => s_locks_lower_in(38,10),
			in1                => s_in1(38,10),
			in2                => s_in2(38,10),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(10)
		);
	s_in1(38,10)            <= s_out1(39,10);
	s_in2(38,10)            <= s_out2(39,11);
	s_locks_lower_in(38,10) <= s_locks_lower_out(39,10);

		normal_cell_38_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,11),
			fetch              => s_fetch(38,11),
			data_in            => s_data_in(38,11),
			data_out           => s_data_out(38,11),
			out1               => s_out1(38,11),
			out2               => s_out2(38,11),
			lock_lower_row_out => s_locks_lower_out(38,11),
			lock_lower_row_in  => s_locks_lower_in(38,11),
			in1                => s_in1(38,11),
			in2                => s_in2(38,11),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(11)
		);
	s_in1(38,11)            <= s_out1(39,11);
	s_in2(38,11)            <= s_out2(39,12);
	s_locks_lower_in(38,11) <= s_locks_lower_out(39,11);

		normal_cell_38_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,12),
			fetch              => s_fetch(38,12),
			data_in            => s_data_in(38,12),
			data_out           => s_data_out(38,12),
			out1               => s_out1(38,12),
			out2               => s_out2(38,12),
			lock_lower_row_out => s_locks_lower_out(38,12),
			lock_lower_row_in  => s_locks_lower_in(38,12),
			in1                => s_in1(38,12),
			in2                => s_in2(38,12),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(12)
		);
	s_in1(38,12)            <= s_out1(39,12);
	s_in2(38,12)            <= s_out2(39,13);
	s_locks_lower_in(38,12) <= s_locks_lower_out(39,12);

		normal_cell_38_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,13),
			fetch              => s_fetch(38,13),
			data_in            => s_data_in(38,13),
			data_out           => s_data_out(38,13),
			out1               => s_out1(38,13),
			out2               => s_out2(38,13),
			lock_lower_row_out => s_locks_lower_out(38,13),
			lock_lower_row_in  => s_locks_lower_in(38,13),
			in1                => s_in1(38,13),
			in2                => s_in2(38,13),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(13)
		);
	s_in1(38,13)            <= s_out1(39,13);
	s_in2(38,13)            <= s_out2(39,14);
	s_locks_lower_in(38,13) <= s_locks_lower_out(39,13);

		normal_cell_38_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,14),
			fetch              => s_fetch(38,14),
			data_in            => s_data_in(38,14),
			data_out           => s_data_out(38,14),
			out1               => s_out1(38,14),
			out2               => s_out2(38,14),
			lock_lower_row_out => s_locks_lower_out(38,14),
			lock_lower_row_in  => s_locks_lower_in(38,14),
			in1                => s_in1(38,14),
			in2                => s_in2(38,14),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(14)
		);
	s_in1(38,14)            <= s_out1(39,14);
	s_in2(38,14)            <= s_out2(39,15);
	s_locks_lower_in(38,14) <= s_locks_lower_out(39,14);

		normal_cell_38_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,15),
			fetch              => s_fetch(38,15),
			data_in            => s_data_in(38,15),
			data_out           => s_data_out(38,15),
			out1               => s_out1(38,15),
			out2               => s_out2(38,15),
			lock_lower_row_out => s_locks_lower_out(38,15),
			lock_lower_row_in  => s_locks_lower_in(38,15),
			in1                => s_in1(38,15),
			in2                => s_in2(38,15),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(15)
		);
	s_in1(38,15)            <= s_out1(39,15);
	s_in2(38,15)            <= s_out2(39,16);
	s_locks_lower_in(38,15) <= s_locks_lower_out(39,15);

		normal_cell_38_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,16),
			fetch              => s_fetch(38,16),
			data_in            => s_data_in(38,16),
			data_out           => s_data_out(38,16),
			out1               => s_out1(38,16),
			out2               => s_out2(38,16),
			lock_lower_row_out => s_locks_lower_out(38,16),
			lock_lower_row_in  => s_locks_lower_in(38,16),
			in1                => s_in1(38,16),
			in2                => s_in2(38,16),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(16)
		);
	s_in1(38,16)            <= s_out1(39,16);
	s_in2(38,16)            <= s_out2(39,17);
	s_locks_lower_in(38,16) <= s_locks_lower_out(39,16);

		normal_cell_38_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,17),
			fetch              => s_fetch(38,17),
			data_in            => s_data_in(38,17),
			data_out           => s_data_out(38,17),
			out1               => s_out1(38,17),
			out2               => s_out2(38,17),
			lock_lower_row_out => s_locks_lower_out(38,17),
			lock_lower_row_in  => s_locks_lower_in(38,17),
			in1                => s_in1(38,17),
			in2                => s_in2(38,17),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(17)
		);
	s_in1(38,17)            <= s_out1(39,17);
	s_in2(38,17)            <= s_out2(39,18);
	s_locks_lower_in(38,17) <= s_locks_lower_out(39,17);

		normal_cell_38_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,18),
			fetch              => s_fetch(38,18),
			data_in            => s_data_in(38,18),
			data_out           => s_data_out(38,18),
			out1               => s_out1(38,18),
			out2               => s_out2(38,18),
			lock_lower_row_out => s_locks_lower_out(38,18),
			lock_lower_row_in  => s_locks_lower_in(38,18),
			in1                => s_in1(38,18),
			in2                => s_in2(38,18),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(18)
		);
	s_in1(38,18)            <= s_out1(39,18);
	s_in2(38,18)            <= s_out2(39,19);
	s_locks_lower_in(38,18) <= s_locks_lower_out(39,18);

		normal_cell_38_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,19),
			fetch              => s_fetch(38,19),
			data_in            => s_data_in(38,19),
			data_out           => s_data_out(38,19),
			out1               => s_out1(38,19),
			out2               => s_out2(38,19),
			lock_lower_row_out => s_locks_lower_out(38,19),
			lock_lower_row_in  => s_locks_lower_in(38,19),
			in1                => s_in1(38,19),
			in2                => s_in2(38,19),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(19)
		);
	s_in1(38,19)            <= s_out1(39,19);
	s_in2(38,19)            <= s_out2(39,20);
	s_locks_lower_in(38,19) <= s_locks_lower_out(39,19);

		normal_cell_38_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,20),
			fetch              => s_fetch(38,20),
			data_in            => s_data_in(38,20),
			data_out           => s_data_out(38,20),
			out1               => s_out1(38,20),
			out2               => s_out2(38,20),
			lock_lower_row_out => s_locks_lower_out(38,20),
			lock_lower_row_in  => s_locks_lower_in(38,20),
			in1                => s_in1(38,20),
			in2                => s_in2(38,20),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(20)
		);
	s_in1(38,20)            <= s_out1(39,20);
	s_in2(38,20)            <= s_out2(39,21);
	s_locks_lower_in(38,20) <= s_locks_lower_out(39,20);

		normal_cell_38_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,21),
			fetch              => s_fetch(38,21),
			data_in            => s_data_in(38,21),
			data_out           => s_data_out(38,21),
			out1               => s_out1(38,21),
			out2               => s_out2(38,21),
			lock_lower_row_out => s_locks_lower_out(38,21),
			lock_lower_row_in  => s_locks_lower_in(38,21),
			in1                => s_in1(38,21),
			in2                => s_in2(38,21),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(21)
		);
	s_in1(38,21)            <= s_out1(39,21);
	s_in2(38,21)            <= s_out2(39,22);
	s_locks_lower_in(38,21) <= s_locks_lower_out(39,21);

		normal_cell_38_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,22),
			fetch              => s_fetch(38,22),
			data_in            => s_data_in(38,22),
			data_out           => s_data_out(38,22),
			out1               => s_out1(38,22),
			out2               => s_out2(38,22),
			lock_lower_row_out => s_locks_lower_out(38,22),
			lock_lower_row_in  => s_locks_lower_in(38,22),
			in1                => s_in1(38,22),
			in2                => s_in2(38,22),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(22)
		);
	s_in1(38,22)            <= s_out1(39,22);
	s_in2(38,22)            <= s_out2(39,23);
	s_locks_lower_in(38,22) <= s_locks_lower_out(39,22);

		normal_cell_38_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,23),
			fetch              => s_fetch(38,23),
			data_in            => s_data_in(38,23),
			data_out           => s_data_out(38,23),
			out1               => s_out1(38,23),
			out2               => s_out2(38,23),
			lock_lower_row_out => s_locks_lower_out(38,23),
			lock_lower_row_in  => s_locks_lower_in(38,23),
			in1                => s_in1(38,23),
			in2                => s_in2(38,23),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(23)
		);
	s_in1(38,23)            <= s_out1(39,23);
	s_in2(38,23)            <= s_out2(39,24);
	s_locks_lower_in(38,23) <= s_locks_lower_out(39,23);

		normal_cell_38_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,24),
			fetch              => s_fetch(38,24),
			data_in            => s_data_in(38,24),
			data_out           => s_data_out(38,24),
			out1               => s_out1(38,24),
			out2               => s_out2(38,24),
			lock_lower_row_out => s_locks_lower_out(38,24),
			lock_lower_row_in  => s_locks_lower_in(38,24),
			in1                => s_in1(38,24),
			in2                => s_in2(38,24),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(24)
		);
	s_in1(38,24)            <= s_out1(39,24);
	s_in2(38,24)            <= s_out2(39,25);
	s_locks_lower_in(38,24) <= s_locks_lower_out(39,24);

		normal_cell_38_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,25),
			fetch              => s_fetch(38,25),
			data_in            => s_data_in(38,25),
			data_out           => s_data_out(38,25),
			out1               => s_out1(38,25),
			out2               => s_out2(38,25),
			lock_lower_row_out => s_locks_lower_out(38,25),
			lock_lower_row_in  => s_locks_lower_in(38,25),
			in1                => s_in1(38,25),
			in2                => s_in2(38,25),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(25)
		);
	s_in1(38,25)            <= s_out1(39,25);
	s_in2(38,25)            <= s_out2(39,26);
	s_locks_lower_in(38,25) <= s_locks_lower_out(39,25);

		normal_cell_38_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,26),
			fetch              => s_fetch(38,26),
			data_in            => s_data_in(38,26),
			data_out           => s_data_out(38,26),
			out1               => s_out1(38,26),
			out2               => s_out2(38,26),
			lock_lower_row_out => s_locks_lower_out(38,26),
			lock_lower_row_in  => s_locks_lower_in(38,26),
			in1                => s_in1(38,26),
			in2                => s_in2(38,26),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(26)
		);
	s_in1(38,26)            <= s_out1(39,26);
	s_in2(38,26)            <= s_out2(39,27);
	s_locks_lower_in(38,26) <= s_locks_lower_out(39,26);

		normal_cell_38_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,27),
			fetch              => s_fetch(38,27),
			data_in            => s_data_in(38,27),
			data_out           => s_data_out(38,27),
			out1               => s_out1(38,27),
			out2               => s_out2(38,27),
			lock_lower_row_out => s_locks_lower_out(38,27),
			lock_lower_row_in  => s_locks_lower_in(38,27),
			in1                => s_in1(38,27),
			in2                => s_in2(38,27),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(27)
		);
	s_in1(38,27)            <= s_out1(39,27);
	s_in2(38,27)            <= s_out2(39,28);
	s_locks_lower_in(38,27) <= s_locks_lower_out(39,27);

		normal_cell_38_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,28),
			fetch              => s_fetch(38,28),
			data_in            => s_data_in(38,28),
			data_out           => s_data_out(38,28),
			out1               => s_out1(38,28),
			out2               => s_out2(38,28),
			lock_lower_row_out => s_locks_lower_out(38,28),
			lock_lower_row_in  => s_locks_lower_in(38,28),
			in1                => s_in1(38,28),
			in2                => s_in2(38,28),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(28)
		);
	s_in1(38,28)            <= s_out1(39,28);
	s_in2(38,28)            <= s_out2(39,29);
	s_locks_lower_in(38,28) <= s_locks_lower_out(39,28);

		normal_cell_38_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,29),
			fetch              => s_fetch(38,29),
			data_in            => s_data_in(38,29),
			data_out           => s_data_out(38,29),
			out1               => s_out1(38,29),
			out2               => s_out2(38,29),
			lock_lower_row_out => s_locks_lower_out(38,29),
			lock_lower_row_in  => s_locks_lower_in(38,29),
			in1                => s_in1(38,29),
			in2                => s_in2(38,29),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(29)
		);
	s_in1(38,29)            <= s_out1(39,29);
	s_in2(38,29)            <= s_out2(39,30);
	s_locks_lower_in(38,29) <= s_locks_lower_out(39,29);

		normal_cell_38_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,30),
			fetch              => s_fetch(38,30),
			data_in            => s_data_in(38,30),
			data_out           => s_data_out(38,30),
			out1               => s_out1(38,30),
			out2               => s_out2(38,30),
			lock_lower_row_out => s_locks_lower_out(38,30),
			lock_lower_row_in  => s_locks_lower_in(38,30),
			in1                => s_in1(38,30),
			in2                => s_in2(38,30),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(30)
		);
	s_in1(38,30)            <= s_out1(39,30);
	s_in2(38,30)            <= s_out2(39,31);
	s_locks_lower_in(38,30) <= s_locks_lower_out(39,30);

		normal_cell_38_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,31),
			fetch              => s_fetch(38,31),
			data_in            => s_data_in(38,31),
			data_out           => s_data_out(38,31),
			out1               => s_out1(38,31),
			out2               => s_out2(38,31),
			lock_lower_row_out => s_locks_lower_out(38,31),
			lock_lower_row_in  => s_locks_lower_in(38,31),
			in1                => s_in1(38,31),
			in2                => s_in2(38,31),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(31)
		);
	s_in1(38,31)            <= s_out1(39,31);
	s_in2(38,31)            <= s_out2(39,32);
	s_locks_lower_in(38,31) <= s_locks_lower_out(39,31);

		normal_cell_38_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,32),
			fetch              => s_fetch(38,32),
			data_in            => s_data_in(38,32),
			data_out           => s_data_out(38,32),
			out1               => s_out1(38,32),
			out2               => s_out2(38,32),
			lock_lower_row_out => s_locks_lower_out(38,32),
			lock_lower_row_in  => s_locks_lower_in(38,32),
			in1                => s_in1(38,32),
			in2                => s_in2(38,32),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(32)
		);
	s_in1(38,32)            <= s_out1(39,32);
	s_in2(38,32)            <= s_out2(39,33);
	s_locks_lower_in(38,32) <= s_locks_lower_out(39,32);

		normal_cell_38_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,33),
			fetch              => s_fetch(38,33),
			data_in            => s_data_in(38,33),
			data_out           => s_data_out(38,33),
			out1               => s_out1(38,33),
			out2               => s_out2(38,33),
			lock_lower_row_out => s_locks_lower_out(38,33),
			lock_lower_row_in  => s_locks_lower_in(38,33),
			in1                => s_in1(38,33),
			in2                => s_in2(38,33),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(33)
		);
	s_in1(38,33)            <= s_out1(39,33);
	s_in2(38,33)            <= s_out2(39,34);
	s_locks_lower_in(38,33) <= s_locks_lower_out(39,33);

		normal_cell_38_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,34),
			fetch              => s_fetch(38,34),
			data_in            => s_data_in(38,34),
			data_out           => s_data_out(38,34),
			out1               => s_out1(38,34),
			out2               => s_out2(38,34),
			lock_lower_row_out => s_locks_lower_out(38,34),
			lock_lower_row_in  => s_locks_lower_in(38,34),
			in1                => s_in1(38,34),
			in2                => s_in2(38,34),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(34)
		);
	s_in1(38,34)            <= s_out1(39,34);
	s_in2(38,34)            <= s_out2(39,35);
	s_locks_lower_in(38,34) <= s_locks_lower_out(39,34);

		normal_cell_38_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,35),
			fetch              => s_fetch(38,35),
			data_in            => s_data_in(38,35),
			data_out           => s_data_out(38,35),
			out1               => s_out1(38,35),
			out2               => s_out2(38,35),
			lock_lower_row_out => s_locks_lower_out(38,35),
			lock_lower_row_in  => s_locks_lower_in(38,35),
			in1                => s_in1(38,35),
			in2                => s_in2(38,35),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(35)
		);
	s_in1(38,35)            <= s_out1(39,35);
	s_in2(38,35)            <= s_out2(39,36);
	s_locks_lower_in(38,35) <= s_locks_lower_out(39,35);

		normal_cell_38_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,36),
			fetch              => s_fetch(38,36),
			data_in            => s_data_in(38,36),
			data_out           => s_data_out(38,36),
			out1               => s_out1(38,36),
			out2               => s_out2(38,36),
			lock_lower_row_out => s_locks_lower_out(38,36),
			lock_lower_row_in  => s_locks_lower_in(38,36),
			in1                => s_in1(38,36),
			in2                => s_in2(38,36),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(36)
		);
	s_in1(38,36)            <= s_out1(39,36);
	s_in2(38,36)            <= s_out2(39,37);
	s_locks_lower_in(38,36) <= s_locks_lower_out(39,36);

		normal_cell_38_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,37),
			fetch              => s_fetch(38,37),
			data_in            => s_data_in(38,37),
			data_out           => s_data_out(38,37),
			out1               => s_out1(38,37),
			out2               => s_out2(38,37),
			lock_lower_row_out => s_locks_lower_out(38,37),
			lock_lower_row_in  => s_locks_lower_in(38,37),
			in1                => s_in1(38,37),
			in2                => s_in2(38,37),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(37)
		);
	s_in1(38,37)            <= s_out1(39,37);
	s_in2(38,37)            <= s_out2(39,38);
	s_locks_lower_in(38,37) <= s_locks_lower_out(39,37);

		normal_cell_38_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,38),
			fetch              => s_fetch(38,38),
			data_in            => s_data_in(38,38),
			data_out           => s_data_out(38,38),
			out1               => s_out1(38,38),
			out2               => s_out2(38,38),
			lock_lower_row_out => s_locks_lower_out(38,38),
			lock_lower_row_in  => s_locks_lower_in(38,38),
			in1                => s_in1(38,38),
			in2                => s_in2(38,38),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(38)
		);
	s_in1(38,38)            <= s_out1(39,38);
	s_in2(38,38)            <= s_out2(39,39);
	s_locks_lower_in(38,38) <= s_locks_lower_out(39,38);

		normal_cell_38_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,39),
			fetch              => s_fetch(38,39),
			data_in            => s_data_in(38,39),
			data_out           => s_data_out(38,39),
			out1               => s_out1(38,39),
			out2               => s_out2(38,39),
			lock_lower_row_out => s_locks_lower_out(38,39),
			lock_lower_row_in  => s_locks_lower_in(38,39),
			in1                => s_in1(38,39),
			in2                => s_in2(38,39),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(39)
		);
	s_in1(38,39)            <= s_out1(39,39);
	s_in2(38,39)            <= s_out2(39,40);
	s_locks_lower_in(38,39) <= s_locks_lower_out(39,39);

		normal_cell_38_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,40),
			fetch              => s_fetch(38,40),
			data_in            => s_data_in(38,40),
			data_out           => s_data_out(38,40),
			out1               => s_out1(38,40),
			out2               => s_out2(38,40),
			lock_lower_row_out => s_locks_lower_out(38,40),
			lock_lower_row_in  => s_locks_lower_in(38,40),
			in1                => s_in1(38,40),
			in2                => s_in2(38,40),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(40)
		);
	s_in1(38,40)            <= s_out1(39,40);
	s_in2(38,40)            <= s_out2(39,41);
	s_locks_lower_in(38,40) <= s_locks_lower_out(39,40);

		normal_cell_38_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,41),
			fetch              => s_fetch(38,41),
			data_in            => s_data_in(38,41),
			data_out           => s_data_out(38,41),
			out1               => s_out1(38,41),
			out2               => s_out2(38,41),
			lock_lower_row_out => s_locks_lower_out(38,41),
			lock_lower_row_in  => s_locks_lower_in(38,41),
			in1                => s_in1(38,41),
			in2                => s_in2(38,41),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(41)
		);
	s_in1(38,41)            <= s_out1(39,41);
	s_in2(38,41)            <= s_out2(39,42);
	s_locks_lower_in(38,41) <= s_locks_lower_out(39,41);

		normal_cell_38_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,42),
			fetch              => s_fetch(38,42),
			data_in            => s_data_in(38,42),
			data_out           => s_data_out(38,42),
			out1               => s_out1(38,42),
			out2               => s_out2(38,42),
			lock_lower_row_out => s_locks_lower_out(38,42),
			lock_lower_row_in  => s_locks_lower_in(38,42),
			in1                => s_in1(38,42),
			in2                => s_in2(38,42),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(42)
		);
	s_in1(38,42)            <= s_out1(39,42);
	s_in2(38,42)            <= s_out2(39,43);
	s_locks_lower_in(38,42) <= s_locks_lower_out(39,42);

		normal_cell_38_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,43),
			fetch              => s_fetch(38,43),
			data_in            => s_data_in(38,43),
			data_out           => s_data_out(38,43),
			out1               => s_out1(38,43),
			out2               => s_out2(38,43),
			lock_lower_row_out => s_locks_lower_out(38,43),
			lock_lower_row_in  => s_locks_lower_in(38,43),
			in1                => s_in1(38,43),
			in2                => s_in2(38,43),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(43)
		);
	s_in1(38,43)            <= s_out1(39,43);
	s_in2(38,43)            <= s_out2(39,44);
	s_locks_lower_in(38,43) <= s_locks_lower_out(39,43);

		normal_cell_38_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,44),
			fetch              => s_fetch(38,44),
			data_in            => s_data_in(38,44),
			data_out           => s_data_out(38,44),
			out1               => s_out1(38,44),
			out2               => s_out2(38,44),
			lock_lower_row_out => s_locks_lower_out(38,44),
			lock_lower_row_in  => s_locks_lower_in(38,44),
			in1                => s_in1(38,44),
			in2                => s_in2(38,44),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(44)
		);
	s_in1(38,44)            <= s_out1(39,44);
	s_in2(38,44)            <= s_out2(39,45);
	s_locks_lower_in(38,44) <= s_locks_lower_out(39,44);

		normal_cell_38_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,45),
			fetch              => s_fetch(38,45),
			data_in            => s_data_in(38,45),
			data_out           => s_data_out(38,45),
			out1               => s_out1(38,45),
			out2               => s_out2(38,45),
			lock_lower_row_out => s_locks_lower_out(38,45),
			lock_lower_row_in  => s_locks_lower_in(38,45),
			in1                => s_in1(38,45),
			in2                => s_in2(38,45),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(45)
		);
	s_in1(38,45)            <= s_out1(39,45);
	s_in2(38,45)            <= s_out2(39,46);
	s_locks_lower_in(38,45) <= s_locks_lower_out(39,45);

		normal_cell_38_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,46),
			fetch              => s_fetch(38,46),
			data_in            => s_data_in(38,46),
			data_out           => s_data_out(38,46),
			out1               => s_out1(38,46),
			out2               => s_out2(38,46),
			lock_lower_row_out => s_locks_lower_out(38,46),
			lock_lower_row_in  => s_locks_lower_in(38,46),
			in1                => s_in1(38,46),
			in2                => s_in2(38,46),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(46)
		);
	s_in1(38,46)            <= s_out1(39,46);
	s_in2(38,46)            <= s_out2(39,47);
	s_locks_lower_in(38,46) <= s_locks_lower_out(39,46);

		normal_cell_38_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,47),
			fetch              => s_fetch(38,47),
			data_in            => s_data_in(38,47),
			data_out           => s_data_out(38,47),
			out1               => s_out1(38,47),
			out2               => s_out2(38,47),
			lock_lower_row_out => s_locks_lower_out(38,47),
			lock_lower_row_in  => s_locks_lower_in(38,47),
			in1                => s_in1(38,47),
			in2                => s_in2(38,47),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(47)
		);
	s_in1(38,47)            <= s_out1(39,47);
	s_in2(38,47)            <= s_out2(39,48);
	s_locks_lower_in(38,47) <= s_locks_lower_out(39,47);

		normal_cell_38_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,48),
			fetch              => s_fetch(38,48),
			data_in            => s_data_in(38,48),
			data_out           => s_data_out(38,48),
			out1               => s_out1(38,48),
			out2               => s_out2(38,48),
			lock_lower_row_out => s_locks_lower_out(38,48),
			lock_lower_row_in  => s_locks_lower_in(38,48),
			in1                => s_in1(38,48),
			in2                => s_in2(38,48),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(48)
		);
	s_in1(38,48)            <= s_out1(39,48);
	s_in2(38,48)            <= s_out2(39,49);
	s_locks_lower_in(38,48) <= s_locks_lower_out(39,48);

		normal_cell_38_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,49),
			fetch              => s_fetch(38,49),
			data_in            => s_data_in(38,49),
			data_out           => s_data_out(38,49),
			out1               => s_out1(38,49),
			out2               => s_out2(38,49),
			lock_lower_row_out => s_locks_lower_out(38,49),
			lock_lower_row_in  => s_locks_lower_in(38,49),
			in1                => s_in1(38,49),
			in2                => s_in2(38,49),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(49)
		);
	s_in1(38,49)            <= s_out1(39,49);
	s_in2(38,49)            <= s_out2(39,50);
	s_locks_lower_in(38,49) <= s_locks_lower_out(39,49);

		normal_cell_38_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,50),
			fetch              => s_fetch(38,50),
			data_in            => s_data_in(38,50),
			data_out           => s_data_out(38,50),
			out1               => s_out1(38,50),
			out2               => s_out2(38,50),
			lock_lower_row_out => s_locks_lower_out(38,50),
			lock_lower_row_in  => s_locks_lower_in(38,50),
			in1                => s_in1(38,50),
			in2                => s_in2(38,50),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(50)
		);
	s_in1(38,50)            <= s_out1(39,50);
	s_in2(38,50)            <= s_out2(39,51);
	s_locks_lower_in(38,50) <= s_locks_lower_out(39,50);

		normal_cell_38_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,51),
			fetch              => s_fetch(38,51),
			data_in            => s_data_in(38,51),
			data_out           => s_data_out(38,51),
			out1               => s_out1(38,51),
			out2               => s_out2(38,51),
			lock_lower_row_out => s_locks_lower_out(38,51),
			lock_lower_row_in  => s_locks_lower_in(38,51),
			in1                => s_in1(38,51),
			in2                => s_in2(38,51),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(51)
		);
	s_in1(38,51)            <= s_out1(39,51);
	s_in2(38,51)            <= s_out2(39,52);
	s_locks_lower_in(38,51) <= s_locks_lower_out(39,51);

		normal_cell_38_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,52),
			fetch              => s_fetch(38,52),
			data_in            => s_data_in(38,52),
			data_out           => s_data_out(38,52),
			out1               => s_out1(38,52),
			out2               => s_out2(38,52),
			lock_lower_row_out => s_locks_lower_out(38,52),
			lock_lower_row_in  => s_locks_lower_in(38,52),
			in1                => s_in1(38,52),
			in2                => s_in2(38,52),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(52)
		);
	s_in1(38,52)            <= s_out1(39,52);
	s_in2(38,52)            <= s_out2(39,53);
	s_locks_lower_in(38,52) <= s_locks_lower_out(39,52);

		normal_cell_38_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,53),
			fetch              => s_fetch(38,53),
			data_in            => s_data_in(38,53),
			data_out           => s_data_out(38,53),
			out1               => s_out1(38,53),
			out2               => s_out2(38,53),
			lock_lower_row_out => s_locks_lower_out(38,53),
			lock_lower_row_in  => s_locks_lower_in(38,53),
			in1                => s_in1(38,53),
			in2                => s_in2(38,53),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(53)
		);
	s_in1(38,53)            <= s_out1(39,53);
	s_in2(38,53)            <= s_out2(39,54);
	s_locks_lower_in(38,53) <= s_locks_lower_out(39,53);

		normal_cell_38_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,54),
			fetch              => s_fetch(38,54),
			data_in            => s_data_in(38,54),
			data_out           => s_data_out(38,54),
			out1               => s_out1(38,54),
			out2               => s_out2(38,54),
			lock_lower_row_out => s_locks_lower_out(38,54),
			lock_lower_row_in  => s_locks_lower_in(38,54),
			in1                => s_in1(38,54),
			in2                => s_in2(38,54),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(54)
		);
	s_in1(38,54)            <= s_out1(39,54);
	s_in2(38,54)            <= s_out2(39,55);
	s_locks_lower_in(38,54) <= s_locks_lower_out(39,54);

		normal_cell_38_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,55),
			fetch              => s_fetch(38,55),
			data_in            => s_data_in(38,55),
			data_out           => s_data_out(38,55),
			out1               => s_out1(38,55),
			out2               => s_out2(38,55),
			lock_lower_row_out => s_locks_lower_out(38,55),
			lock_lower_row_in  => s_locks_lower_in(38,55),
			in1                => s_in1(38,55),
			in2                => s_in2(38,55),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(55)
		);
	s_in1(38,55)            <= s_out1(39,55);
	s_in2(38,55)            <= s_out2(39,56);
	s_locks_lower_in(38,55) <= s_locks_lower_out(39,55);

		normal_cell_38_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,56),
			fetch              => s_fetch(38,56),
			data_in            => s_data_in(38,56),
			data_out           => s_data_out(38,56),
			out1               => s_out1(38,56),
			out2               => s_out2(38,56),
			lock_lower_row_out => s_locks_lower_out(38,56),
			lock_lower_row_in  => s_locks_lower_in(38,56),
			in1                => s_in1(38,56),
			in2                => s_in2(38,56),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(56)
		);
	s_in1(38,56)            <= s_out1(39,56);
	s_in2(38,56)            <= s_out2(39,57);
	s_locks_lower_in(38,56) <= s_locks_lower_out(39,56);

		normal_cell_38_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,57),
			fetch              => s_fetch(38,57),
			data_in            => s_data_in(38,57),
			data_out           => s_data_out(38,57),
			out1               => s_out1(38,57),
			out2               => s_out2(38,57),
			lock_lower_row_out => s_locks_lower_out(38,57),
			lock_lower_row_in  => s_locks_lower_in(38,57),
			in1                => s_in1(38,57),
			in2                => s_in2(38,57),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(57)
		);
	s_in1(38,57)            <= s_out1(39,57);
	s_in2(38,57)            <= s_out2(39,58);
	s_locks_lower_in(38,57) <= s_locks_lower_out(39,57);

		normal_cell_38_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,58),
			fetch              => s_fetch(38,58),
			data_in            => s_data_in(38,58),
			data_out           => s_data_out(38,58),
			out1               => s_out1(38,58),
			out2               => s_out2(38,58),
			lock_lower_row_out => s_locks_lower_out(38,58),
			lock_lower_row_in  => s_locks_lower_in(38,58),
			in1                => s_in1(38,58),
			in2                => s_in2(38,58),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(58)
		);
	s_in1(38,58)            <= s_out1(39,58);
	s_in2(38,58)            <= s_out2(39,59);
	s_locks_lower_in(38,58) <= s_locks_lower_out(39,58);

		normal_cell_38_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,59),
			fetch              => s_fetch(38,59),
			data_in            => s_data_in(38,59),
			data_out           => s_data_out(38,59),
			out1               => s_out1(38,59),
			out2               => s_out2(38,59),
			lock_lower_row_out => s_locks_lower_out(38,59),
			lock_lower_row_in  => s_locks_lower_in(38,59),
			in1                => s_in1(38,59),
			in2                => s_in2(38,59),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(59)
		);
	s_in1(38,59)            <= s_out1(39,59);
	s_in2(38,59)            <= s_out2(39,60);
	s_locks_lower_in(38,59) <= s_locks_lower_out(39,59);

		last_col_cell_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(38,60),
			fetch              => s_fetch(38,60),
			data_in            => s_data_in(38,60),
			data_out           => s_data_out(38,60),
			out1               => s_out1(38,60),
			out2               => s_out2(38,60),
			lock_lower_row_out => s_locks_lower_out(38,60),
			lock_lower_row_in  => s_locks_lower_in(38,60),
			in1                => s_in1(38,60),
			in2                => (others => '0'),
			lock_row           => s_locks(38),
			piv_found          => s_piv_found,
			row_data           => s_row_data(38),
			col_data           => s_col_data(60)
		);
	s_in1(38,60)            <= s_out1(39,60);
	s_locks_lower_in(38,60) <= s_locks_lower_out(39,60);

		normal_cell_39_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,1),
			fetch              => s_fetch(39,1),
			data_in            => s_data_in(39,1),
			data_out           => s_data_out(39,1),
			out1               => s_out1(39,1),
			out2               => s_out2(39,1),
			lock_lower_row_out => s_locks_lower_out(39,1),
			lock_lower_row_in  => s_locks_lower_in(39,1),
			in1                => s_in1(39,1),
			in2                => s_in2(39,1),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(1)
		);
	s_in1(39,1)            <= s_out1(40,1);
	s_in2(39,1)            <= s_out2(40,2);
	s_locks_lower_in(39,1) <= s_locks_lower_out(40,1);

		normal_cell_39_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,2),
			fetch              => s_fetch(39,2),
			data_in            => s_data_in(39,2),
			data_out           => s_data_out(39,2),
			out1               => s_out1(39,2),
			out2               => s_out2(39,2),
			lock_lower_row_out => s_locks_lower_out(39,2),
			lock_lower_row_in  => s_locks_lower_in(39,2),
			in1                => s_in1(39,2),
			in2                => s_in2(39,2),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(2)
		);
	s_in1(39,2)            <= s_out1(40,2);
	s_in2(39,2)            <= s_out2(40,3);
	s_locks_lower_in(39,2) <= s_locks_lower_out(40,2);

		normal_cell_39_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,3),
			fetch              => s_fetch(39,3),
			data_in            => s_data_in(39,3),
			data_out           => s_data_out(39,3),
			out1               => s_out1(39,3),
			out2               => s_out2(39,3),
			lock_lower_row_out => s_locks_lower_out(39,3),
			lock_lower_row_in  => s_locks_lower_in(39,3),
			in1                => s_in1(39,3),
			in2                => s_in2(39,3),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(3)
		);
	s_in1(39,3)            <= s_out1(40,3);
	s_in2(39,3)            <= s_out2(40,4);
	s_locks_lower_in(39,3) <= s_locks_lower_out(40,3);

		normal_cell_39_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,4),
			fetch              => s_fetch(39,4),
			data_in            => s_data_in(39,4),
			data_out           => s_data_out(39,4),
			out1               => s_out1(39,4),
			out2               => s_out2(39,4),
			lock_lower_row_out => s_locks_lower_out(39,4),
			lock_lower_row_in  => s_locks_lower_in(39,4),
			in1                => s_in1(39,4),
			in2                => s_in2(39,4),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(4)
		);
	s_in1(39,4)            <= s_out1(40,4);
	s_in2(39,4)            <= s_out2(40,5);
	s_locks_lower_in(39,4) <= s_locks_lower_out(40,4);

		normal_cell_39_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,5),
			fetch              => s_fetch(39,5),
			data_in            => s_data_in(39,5),
			data_out           => s_data_out(39,5),
			out1               => s_out1(39,5),
			out2               => s_out2(39,5),
			lock_lower_row_out => s_locks_lower_out(39,5),
			lock_lower_row_in  => s_locks_lower_in(39,5),
			in1                => s_in1(39,5),
			in2                => s_in2(39,5),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(5)
		);
	s_in1(39,5)            <= s_out1(40,5);
	s_in2(39,5)            <= s_out2(40,6);
	s_locks_lower_in(39,5) <= s_locks_lower_out(40,5);

		normal_cell_39_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,6),
			fetch              => s_fetch(39,6),
			data_in            => s_data_in(39,6),
			data_out           => s_data_out(39,6),
			out1               => s_out1(39,6),
			out2               => s_out2(39,6),
			lock_lower_row_out => s_locks_lower_out(39,6),
			lock_lower_row_in  => s_locks_lower_in(39,6),
			in1                => s_in1(39,6),
			in2                => s_in2(39,6),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(6)
		);
	s_in1(39,6)            <= s_out1(40,6);
	s_in2(39,6)            <= s_out2(40,7);
	s_locks_lower_in(39,6) <= s_locks_lower_out(40,6);

		normal_cell_39_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,7),
			fetch              => s_fetch(39,7),
			data_in            => s_data_in(39,7),
			data_out           => s_data_out(39,7),
			out1               => s_out1(39,7),
			out2               => s_out2(39,7),
			lock_lower_row_out => s_locks_lower_out(39,7),
			lock_lower_row_in  => s_locks_lower_in(39,7),
			in1                => s_in1(39,7),
			in2                => s_in2(39,7),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(7)
		);
	s_in1(39,7)            <= s_out1(40,7);
	s_in2(39,7)            <= s_out2(40,8);
	s_locks_lower_in(39,7) <= s_locks_lower_out(40,7);

		normal_cell_39_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,8),
			fetch              => s_fetch(39,8),
			data_in            => s_data_in(39,8),
			data_out           => s_data_out(39,8),
			out1               => s_out1(39,8),
			out2               => s_out2(39,8),
			lock_lower_row_out => s_locks_lower_out(39,8),
			lock_lower_row_in  => s_locks_lower_in(39,8),
			in1                => s_in1(39,8),
			in2                => s_in2(39,8),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(8)
		);
	s_in1(39,8)            <= s_out1(40,8);
	s_in2(39,8)            <= s_out2(40,9);
	s_locks_lower_in(39,8) <= s_locks_lower_out(40,8);

		normal_cell_39_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,9),
			fetch              => s_fetch(39,9),
			data_in            => s_data_in(39,9),
			data_out           => s_data_out(39,9),
			out1               => s_out1(39,9),
			out2               => s_out2(39,9),
			lock_lower_row_out => s_locks_lower_out(39,9),
			lock_lower_row_in  => s_locks_lower_in(39,9),
			in1                => s_in1(39,9),
			in2                => s_in2(39,9),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(9)
		);
	s_in1(39,9)            <= s_out1(40,9);
	s_in2(39,9)            <= s_out2(40,10);
	s_locks_lower_in(39,9) <= s_locks_lower_out(40,9);

		normal_cell_39_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,10),
			fetch              => s_fetch(39,10),
			data_in            => s_data_in(39,10),
			data_out           => s_data_out(39,10),
			out1               => s_out1(39,10),
			out2               => s_out2(39,10),
			lock_lower_row_out => s_locks_lower_out(39,10),
			lock_lower_row_in  => s_locks_lower_in(39,10),
			in1                => s_in1(39,10),
			in2                => s_in2(39,10),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(10)
		);
	s_in1(39,10)            <= s_out1(40,10);
	s_in2(39,10)            <= s_out2(40,11);
	s_locks_lower_in(39,10) <= s_locks_lower_out(40,10);

		normal_cell_39_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,11),
			fetch              => s_fetch(39,11),
			data_in            => s_data_in(39,11),
			data_out           => s_data_out(39,11),
			out1               => s_out1(39,11),
			out2               => s_out2(39,11),
			lock_lower_row_out => s_locks_lower_out(39,11),
			lock_lower_row_in  => s_locks_lower_in(39,11),
			in1                => s_in1(39,11),
			in2                => s_in2(39,11),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(11)
		);
	s_in1(39,11)            <= s_out1(40,11);
	s_in2(39,11)            <= s_out2(40,12);
	s_locks_lower_in(39,11) <= s_locks_lower_out(40,11);

		normal_cell_39_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,12),
			fetch              => s_fetch(39,12),
			data_in            => s_data_in(39,12),
			data_out           => s_data_out(39,12),
			out1               => s_out1(39,12),
			out2               => s_out2(39,12),
			lock_lower_row_out => s_locks_lower_out(39,12),
			lock_lower_row_in  => s_locks_lower_in(39,12),
			in1                => s_in1(39,12),
			in2                => s_in2(39,12),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(12)
		);
	s_in1(39,12)            <= s_out1(40,12);
	s_in2(39,12)            <= s_out2(40,13);
	s_locks_lower_in(39,12) <= s_locks_lower_out(40,12);

		normal_cell_39_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,13),
			fetch              => s_fetch(39,13),
			data_in            => s_data_in(39,13),
			data_out           => s_data_out(39,13),
			out1               => s_out1(39,13),
			out2               => s_out2(39,13),
			lock_lower_row_out => s_locks_lower_out(39,13),
			lock_lower_row_in  => s_locks_lower_in(39,13),
			in1                => s_in1(39,13),
			in2                => s_in2(39,13),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(13)
		);
	s_in1(39,13)            <= s_out1(40,13);
	s_in2(39,13)            <= s_out2(40,14);
	s_locks_lower_in(39,13) <= s_locks_lower_out(40,13);

		normal_cell_39_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,14),
			fetch              => s_fetch(39,14),
			data_in            => s_data_in(39,14),
			data_out           => s_data_out(39,14),
			out1               => s_out1(39,14),
			out2               => s_out2(39,14),
			lock_lower_row_out => s_locks_lower_out(39,14),
			lock_lower_row_in  => s_locks_lower_in(39,14),
			in1                => s_in1(39,14),
			in2                => s_in2(39,14),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(14)
		);
	s_in1(39,14)            <= s_out1(40,14);
	s_in2(39,14)            <= s_out2(40,15);
	s_locks_lower_in(39,14) <= s_locks_lower_out(40,14);

		normal_cell_39_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,15),
			fetch              => s_fetch(39,15),
			data_in            => s_data_in(39,15),
			data_out           => s_data_out(39,15),
			out1               => s_out1(39,15),
			out2               => s_out2(39,15),
			lock_lower_row_out => s_locks_lower_out(39,15),
			lock_lower_row_in  => s_locks_lower_in(39,15),
			in1                => s_in1(39,15),
			in2                => s_in2(39,15),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(15)
		);
	s_in1(39,15)            <= s_out1(40,15);
	s_in2(39,15)            <= s_out2(40,16);
	s_locks_lower_in(39,15) <= s_locks_lower_out(40,15);

		normal_cell_39_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,16),
			fetch              => s_fetch(39,16),
			data_in            => s_data_in(39,16),
			data_out           => s_data_out(39,16),
			out1               => s_out1(39,16),
			out2               => s_out2(39,16),
			lock_lower_row_out => s_locks_lower_out(39,16),
			lock_lower_row_in  => s_locks_lower_in(39,16),
			in1                => s_in1(39,16),
			in2                => s_in2(39,16),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(16)
		);
	s_in1(39,16)            <= s_out1(40,16);
	s_in2(39,16)            <= s_out2(40,17);
	s_locks_lower_in(39,16) <= s_locks_lower_out(40,16);

		normal_cell_39_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,17),
			fetch              => s_fetch(39,17),
			data_in            => s_data_in(39,17),
			data_out           => s_data_out(39,17),
			out1               => s_out1(39,17),
			out2               => s_out2(39,17),
			lock_lower_row_out => s_locks_lower_out(39,17),
			lock_lower_row_in  => s_locks_lower_in(39,17),
			in1                => s_in1(39,17),
			in2                => s_in2(39,17),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(17)
		);
	s_in1(39,17)            <= s_out1(40,17);
	s_in2(39,17)            <= s_out2(40,18);
	s_locks_lower_in(39,17) <= s_locks_lower_out(40,17);

		normal_cell_39_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,18),
			fetch              => s_fetch(39,18),
			data_in            => s_data_in(39,18),
			data_out           => s_data_out(39,18),
			out1               => s_out1(39,18),
			out2               => s_out2(39,18),
			lock_lower_row_out => s_locks_lower_out(39,18),
			lock_lower_row_in  => s_locks_lower_in(39,18),
			in1                => s_in1(39,18),
			in2                => s_in2(39,18),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(18)
		);
	s_in1(39,18)            <= s_out1(40,18);
	s_in2(39,18)            <= s_out2(40,19);
	s_locks_lower_in(39,18) <= s_locks_lower_out(40,18);

		normal_cell_39_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,19),
			fetch              => s_fetch(39,19),
			data_in            => s_data_in(39,19),
			data_out           => s_data_out(39,19),
			out1               => s_out1(39,19),
			out2               => s_out2(39,19),
			lock_lower_row_out => s_locks_lower_out(39,19),
			lock_lower_row_in  => s_locks_lower_in(39,19),
			in1                => s_in1(39,19),
			in2                => s_in2(39,19),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(19)
		);
	s_in1(39,19)            <= s_out1(40,19);
	s_in2(39,19)            <= s_out2(40,20);
	s_locks_lower_in(39,19) <= s_locks_lower_out(40,19);

		normal_cell_39_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,20),
			fetch              => s_fetch(39,20),
			data_in            => s_data_in(39,20),
			data_out           => s_data_out(39,20),
			out1               => s_out1(39,20),
			out2               => s_out2(39,20),
			lock_lower_row_out => s_locks_lower_out(39,20),
			lock_lower_row_in  => s_locks_lower_in(39,20),
			in1                => s_in1(39,20),
			in2                => s_in2(39,20),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(20)
		);
	s_in1(39,20)            <= s_out1(40,20);
	s_in2(39,20)            <= s_out2(40,21);
	s_locks_lower_in(39,20) <= s_locks_lower_out(40,20);

		normal_cell_39_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,21),
			fetch              => s_fetch(39,21),
			data_in            => s_data_in(39,21),
			data_out           => s_data_out(39,21),
			out1               => s_out1(39,21),
			out2               => s_out2(39,21),
			lock_lower_row_out => s_locks_lower_out(39,21),
			lock_lower_row_in  => s_locks_lower_in(39,21),
			in1                => s_in1(39,21),
			in2                => s_in2(39,21),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(21)
		);
	s_in1(39,21)            <= s_out1(40,21);
	s_in2(39,21)            <= s_out2(40,22);
	s_locks_lower_in(39,21) <= s_locks_lower_out(40,21);

		normal_cell_39_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,22),
			fetch              => s_fetch(39,22),
			data_in            => s_data_in(39,22),
			data_out           => s_data_out(39,22),
			out1               => s_out1(39,22),
			out2               => s_out2(39,22),
			lock_lower_row_out => s_locks_lower_out(39,22),
			lock_lower_row_in  => s_locks_lower_in(39,22),
			in1                => s_in1(39,22),
			in2                => s_in2(39,22),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(22)
		);
	s_in1(39,22)            <= s_out1(40,22);
	s_in2(39,22)            <= s_out2(40,23);
	s_locks_lower_in(39,22) <= s_locks_lower_out(40,22);

		normal_cell_39_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,23),
			fetch              => s_fetch(39,23),
			data_in            => s_data_in(39,23),
			data_out           => s_data_out(39,23),
			out1               => s_out1(39,23),
			out2               => s_out2(39,23),
			lock_lower_row_out => s_locks_lower_out(39,23),
			lock_lower_row_in  => s_locks_lower_in(39,23),
			in1                => s_in1(39,23),
			in2                => s_in2(39,23),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(23)
		);
	s_in1(39,23)            <= s_out1(40,23);
	s_in2(39,23)            <= s_out2(40,24);
	s_locks_lower_in(39,23) <= s_locks_lower_out(40,23);

		normal_cell_39_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,24),
			fetch              => s_fetch(39,24),
			data_in            => s_data_in(39,24),
			data_out           => s_data_out(39,24),
			out1               => s_out1(39,24),
			out2               => s_out2(39,24),
			lock_lower_row_out => s_locks_lower_out(39,24),
			lock_lower_row_in  => s_locks_lower_in(39,24),
			in1                => s_in1(39,24),
			in2                => s_in2(39,24),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(24)
		);
	s_in1(39,24)            <= s_out1(40,24);
	s_in2(39,24)            <= s_out2(40,25);
	s_locks_lower_in(39,24) <= s_locks_lower_out(40,24);

		normal_cell_39_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,25),
			fetch              => s_fetch(39,25),
			data_in            => s_data_in(39,25),
			data_out           => s_data_out(39,25),
			out1               => s_out1(39,25),
			out2               => s_out2(39,25),
			lock_lower_row_out => s_locks_lower_out(39,25),
			lock_lower_row_in  => s_locks_lower_in(39,25),
			in1                => s_in1(39,25),
			in2                => s_in2(39,25),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(25)
		);
	s_in1(39,25)            <= s_out1(40,25);
	s_in2(39,25)            <= s_out2(40,26);
	s_locks_lower_in(39,25) <= s_locks_lower_out(40,25);

		normal_cell_39_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,26),
			fetch              => s_fetch(39,26),
			data_in            => s_data_in(39,26),
			data_out           => s_data_out(39,26),
			out1               => s_out1(39,26),
			out2               => s_out2(39,26),
			lock_lower_row_out => s_locks_lower_out(39,26),
			lock_lower_row_in  => s_locks_lower_in(39,26),
			in1                => s_in1(39,26),
			in2                => s_in2(39,26),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(26)
		);
	s_in1(39,26)            <= s_out1(40,26);
	s_in2(39,26)            <= s_out2(40,27);
	s_locks_lower_in(39,26) <= s_locks_lower_out(40,26);

		normal_cell_39_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,27),
			fetch              => s_fetch(39,27),
			data_in            => s_data_in(39,27),
			data_out           => s_data_out(39,27),
			out1               => s_out1(39,27),
			out2               => s_out2(39,27),
			lock_lower_row_out => s_locks_lower_out(39,27),
			lock_lower_row_in  => s_locks_lower_in(39,27),
			in1                => s_in1(39,27),
			in2                => s_in2(39,27),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(27)
		);
	s_in1(39,27)            <= s_out1(40,27);
	s_in2(39,27)            <= s_out2(40,28);
	s_locks_lower_in(39,27) <= s_locks_lower_out(40,27);

		normal_cell_39_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,28),
			fetch              => s_fetch(39,28),
			data_in            => s_data_in(39,28),
			data_out           => s_data_out(39,28),
			out1               => s_out1(39,28),
			out2               => s_out2(39,28),
			lock_lower_row_out => s_locks_lower_out(39,28),
			lock_lower_row_in  => s_locks_lower_in(39,28),
			in1                => s_in1(39,28),
			in2                => s_in2(39,28),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(28)
		);
	s_in1(39,28)            <= s_out1(40,28);
	s_in2(39,28)            <= s_out2(40,29);
	s_locks_lower_in(39,28) <= s_locks_lower_out(40,28);

		normal_cell_39_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,29),
			fetch              => s_fetch(39,29),
			data_in            => s_data_in(39,29),
			data_out           => s_data_out(39,29),
			out1               => s_out1(39,29),
			out2               => s_out2(39,29),
			lock_lower_row_out => s_locks_lower_out(39,29),
			lock_lower_row_in  => s_locks_lower_in(39,29),
			in1                => s_in1(39,29),
			in2                => s_in2(39,29),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(29)
		);
	s_in1(39,29)            <= s_out1(40,29);
	s_in2(39,29)            <= s_out2(40,30);
	s_locks_lower_in(39,29) <= s_locks_lower_out(40,29);

		normal_cell_39_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,30),
			fetch              => s_fetch(39,30),
			data_in            => s_data_in(39,30),
			data_out           => s_data_out(39,30),
			out1               => s_out1(39,30),
			out2               => s_out2(39,30),
			lock_lower_row_out => s_locks_lower_out(39,30),
			lock_lower_row_in  => s_locks_lower_in(39,30),
			in1                => s_in1(39,30),
			in2                => s_in2(39,30),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(30)
		);
	s_in1(39,30)            <= s_out1(40,30);
	s_in2(39,30)            <= s_out2(40,31);
	s_locks_lower_in(39,30) <= s_locks_lower_out(40,30);

		normal_cell_39_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,31),
			fetch              => s_fetch(39,31),
			data_in            => s_data_in(39,31),
			data_out           => s_data_out(39,31),
			out1               => s_out1(39,31),
			out2               => s_out2(39,31),
			lock_lower_row_out => s_locks_lower_out(39,31),
			lock_lower_row_in  => s_locks_lower_in(39,31),
			in1                => s_in1(39,31),
			in2                => s_in2(39,31),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(31)
		);
	s_in1(39,31)            <= s_out1(40,31);
	s_in2(39,31)            <= s_out2(40,32);
	s_locks_lower_in(39,31) <= s_locks_lower_out(40,31);

		normal_cell_39_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,32),
			fetch              => s_fetch(39,32),
			data_in            => s_data_in(39,32),
			data_out           => s_data_out(39,32),
			out1               => s_out1(39,32),
			out2               => s_out2(39,32),
			lock_lower_row_out => s_locks_lower_out(39,32),
			lock_lower_row_in  => s_locks_lower_in(39,32),
			in1                => s_in1(39,32),
			in2                => s_in2(39,32),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(32)
		);
	s_in1(39,32)            <= s_out1(40,32);
	s_in2(39,32)            <= s_out2(40,33);
	s_locks_lower_in(39,32) <= s_locks_lower_out(40,32);

		normal_cell_39_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,33),
			fetch              => s_fetch(39,33),
			data_in            => s_data_in(39,33),
			data_out           => s_data_out(39,33),
			out1               => s_out1(39,33),
			out2               => s_out2(39,33),
			lock_lower_row_out => s_locks_lower_out(39,33),
			lock_lower_row_in  => s_locks_lower_in(39,33),
			in1                => s_in1(39,33),
			in2                => s_in2(39,33),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(33)
		);
	s_in1(39,33)            <= s_out1(40,33);
	s_in2(39,33)            <= s_out2(40,34);
	s_locks_lower_in(39,33) <= s_locks_lower_out(40,33);

		normal_cell_39_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,34),
			fetch              => s_fetch(39,34),
			data_in            => s_data_in(39,34),
			data_out           => s_data_out(39,34),
			out1               => s_out1(39,34),
			out2               => s_out2(39,34),
			lock_lower_row_out => s_locks_lower_out(39,34),
			lock_lower_row_in  => s_locks_lower_in(39,34),
			in1                => s_in1(39,34),
			in2                => s_in2(39,34),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(34)
		);
	s_in1(39,34)            <= s_out1(40,34);
	s_in2(39,34)            <= s_out2(40,35);
	s_locks_lower_in(39,34) <= s_locks_lower_out(40,34);

		normal_cell_39_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,35),
			fetch              => s_fetch(39,35),
			data_in            => s_data_in(39,35),
			data_out           => s_data_out(39,35),
			out1               => s_out1(39,35),
			out2               => s_out2(39,35),
			lock_lower_row_out => s_locks_lower_out(39,35),
			lock_lower_row_in  => s_locks_lower_in(39,35),
			in1                => s_in1(39,35),
			in2                => s_in2(39,35),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(35)
		);
	s_in1(39,35)            <= s_out1(40,35);
	s_in2(39,35)            <= s_out2(40,36);
	s_locks_lower_in(39,35) <= s_locks_lower_out(40,35);

		normal_cell_39_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,36),
			fetch              => s_fetch(39,36),
			data_in            => s_data_in(39,36),
			data_out           => s_data_out(39,36),
			out1               => s_out1(39,36),
			out2               => s_out2(39,36),
			lock_lower_row_out => s_locks_lower_out(39,36),
			lock_lower_row_in  => s_locks_lower_in(39,36),
			in1                => s_in1(39,36),
			in2                => s_in2(39,36),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(36)
		);
	s_in1(39,36)            <= s_out1(40,36);
	s_in2(39,36)            <= s_out2(40,37);
	s_locks_lower_in(39,36) <= s_locks_lower_out(40,36);

		normal_cell_39_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,37),
			fetch              => s_fetch(39,37),
			data_in            => s_data_in(39,37),
			data_out           => s_data_out(39,37),
			out1               => s_out1(39,37),
			out2               => s_out2(39,37),
			lock_lower_row_out => s_locks_lower_out(39,37),
			lock_lower_row_in  => s_locks_lower_in(39,37),
			in1                => s_in1(39,37),
			in2                => s_in2(39,37),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(37)
		);
	s_in1(39,37)            <= s_out1(40,37);
	s_in2(39,37)            <= s_out2(40,38);
	s_locks_lower_in(39,37) <= s_locks_lower_out(40,37);

		normal_cell_39_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,38),
			fetch              => s_fetch(39,38),
			data_in            => s_data_in(39,38),
			data_out           => s_data_out(39,38),
			out1               => s_out1(39,38),
			out2               => s_out2(39,38),
			lock_lower_row_out => s_locks_lower_out(39,38),
			lock_lower_row_in  => s_locks_lower_in(39,38),
			in1                => s_in1(39,38),
			in2                => s_in2(39,38),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(38)
		);
	s_in1(39,38)            <= s_out1(40,38);
	s_in2(39,38)            <= s_out2(40,39);
	s_locks_lower_in(39,38) <= s_locks_lower_out(40,38);

		normal_cell_39_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,39),
			fetch              => s_fetch(39,39),
			data_in            => s_data_in(39,39),
			data_out           => s_data_out(39,39),
			out1               => s_out1(39,39),
			out2               => s_out2(39,39),
			lock_lower_row_out => s_locks_lower_out(39,39),
			lock_lower_row_in  => s_locks_lower_in(39,39),
			in1                => s_in1(39,39),
			in2                => s_in2(39,39),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(39)
		);
	s_in1(39,39)            <= s_out1(40,39);
	s_in2(39,39)            <= s_out2(40,40);
	s_locks_lower_in(39,39) <= s_locks_lower_out(40,39);

		normal_cell_39_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,40),
			fetch              => s_fetch(39,40),
			data_in            => s_data_in(39,40),
			data_out           => s_data_out(39,40),
			out1               => s_out1(39,40),
			out2               => s_out2(39,40),
			lock_lower_row_out => s_locks_lower_out(39,40),
			lock_lower_row_in  => s_locks_lower_in(39,40),
			in1                => s_in1(39,40),
			in2                => s_in2(39,40),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(40)
		);
	s_in1(39,40)            <= s_out1(40,40);
	s_in2(39,40)            <= s_out2(40,41);
	s_locks_lower_in(39,40) <= s_locks_lower_out(40,40);

		normal_cell_39_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,41),
			fetch              => s_fetch(39,41),
			data_in            => s_data_in(39,41),
			data_out           => s_data_out(39,41),
			out1               => s_out1(39,41),
			out2               => s_out2(39,41),
			lock_lower_row_out => s_locks_lower_out(39,41),
			lock_lower_row_in  => s_locks_lower_in(39,41),
			in1                => s_in1(39,41),
			in2                => s_in2(39,41),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(41)
		);
	s_in1(39,41)            <= s_out1(40,41);
	s_in2(39,41)            <= s_out2(40,42);
	s_locks_lower_in(39,41) <= s_locks_lower_out(40,41);

		normal_cell_39_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,42),
			fetch              => s_fetch(39,42),
			data_in            => s_data_in(39,42),
			data_out           => s_data_out(39,42),
			out1               => s_out1(39,42),
			out2               => s_out2(39,42),
			lock_lower_row_out => s_locks_lower_out(39,42),
			lock_lower_row_in  => s_locks_lower_in(39,42),
			in1                => s_in1(39,42),
			in2                => s_in2(39,42),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(42)
		);
	s_in1(39,42)            <= s_out1(40,42);
	s_in2(39,42)            <= s_out2(40,43);
	s_locks_lower_in(39,42) <= s_locks_lower_out(40,42);

		normal_cell_39_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,43),
			fetch              => s_fetch(39,43),
			data_in            => s_data_in(39,43),
			data_out           => s_data_out(39,43),
			out1               => s_out1(39,43),
			out2               => s_out2(39,43),
			lock_lower_row_out => s_locks_lower_out(39,43),
			lock_lower_row_in  => s_locks_lower_in(39,43),
			in1                => s_in1(39,43),
			in2                => s_in2(39,43),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(43)
		);
	s_in1(39,43)            <= s_out1(40,43);
	s_in2(39,43)            <= s_out2(40,44);
	s_locks_lower_in(39,43) <= s_locks_lower_out(40,43);

		normal_cell_39_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,44),
			fetch              => s_fetch(39,44),
			data_in            => s_data_in(39,44),
			data_out           => s_data_out(39,44),
			out1               => s_out1(39,44),
			out2               => s_out2(39,44),
			lock_lower_row_out => s_locks_lower_out(39,44),
			lock_lower_row_in  => s_locks_lower_in(39,44),
			in1                => s_in1(39,44),
			in2                => s_in2(39,44),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(44)
		);
	s_in1(39,44)            <= s_out1(40,44);
	s_in2(39,44)            <= s_out2(40,45);
	s_locks_lower_in(39,44) <= s_locks_lower_out(40,44);

		normal_cell_39_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,45),
			fetch              => s_fetch(39,45),
			data_in            => s_data_in(39,45),
			data_out           => s_data_out(39,45),
			out1               => s_out1(39,45),
			out2               => s_out2(39,45),
			lock_lower_row_out => s_locks_lower_out(39,45),
			lock_lower_row_in  => s_locks_lower_in(39,45),
			in1                => s_in1(39,45),
			in2                => s_in2(39,45),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(45)
		);
	s_in1(39,45)            <= s_out1(40,45);
	s_in2(39,45)            <= s_out2(40,46);
	s_locks_lower_in(39,45) <= s_locks_lower_out(40,45);

		normal_cell_39_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,46),
			fetch              => s_fetch(39,46),
			data_in            => s_data_in(39,46),
			data_out           => s_data_out(39,46),
			out1               => s_out1(39,46),
			out2               => s_out2(39,46),
			lock_lower_row_out => s_locks_lower_out(39,46),
			lock_lower_row_in  => s_locks_lower_in(39,46),
			in1                => s_in1(39,46),
			in2                => s_in2(39,46),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(46)
		);
	s_in1(39,46)            <= s_out1(40,46);
	s_in2(39,46)            <= s_out2(40,47);
	s_locks_lower_in(39,46) <= s_locks_lower_out(40,46);

		normal_cell_39_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,47),
			fetch              => s_fetch(39,47),
			data_in            => s_data_in(39,47),
			data_out           => s_data_out(39,47),
			out1               => s_out1(39,47),
			out2               => s_out2(39,47),
			lock_lower_row_out => s_locks_lower_out(39,47),
			lock_lower_row_in  => s_locks_lower_in(39,47),
			in1                => s_in1(39,47),
			in2                => s_in2(39,47),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(47)
		);
	s_in1(39,47)            <= s_out1(40,47);
	s_in2(39,47)            <= s_out2(40,48);
	s_locks_lower_in(39,47) <= s_locks_lower_out(40,47);

		normal_cell_39_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,48),
			fetch              => s_fetch(39,48),
			data_in            => s_data_in(39,48),
			data_out           => s_data_out(39,48),
			out1               => s_out1(39,48),
			out2               => s_out2(39,48),
			lock_lower_row_out => s_locks_lower_out(39,48),
			lock_lower_row_in  => s_locks_lower_in(39,48),
			in1                => s_in1(39,48),
			in2                => s_in2(39,48),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(48)
		);
	s_in1(39,48)            <= s_out1(40,48);
	s_in2(39,48)            <= s_out2(40,49);
	s_locks_lower_in(39,48) <= s_locks_lower_out(40,48);

		normal_cell_39_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,49),
			fetch              => s_fetch(39,49),
			data_in            => s_data_in(39,49),
			data_out           => s_data_out(39,49),
			out1               => s_out1(39,49),
			out2               => s_out2(39,49),
			lock_lower_row_out => s_locks_lower_out(39,49),
			lock_lower_row_in  => s_locks_lower_in(39,49),
			in1                => s_in1(39,49),
			in2                => s_in2(39,49),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(49)
		);
	s_in1(39,49)            <= s_out1(40,49);
	s_in2(39,49)            <= s_out2(40,50);
	s_locks_lower_in(39,49) <= s_locks_lower_out(40,49);

		normal_cell_39_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,50),
			fetch              => s_fetch(39,50),
			data_in            => s_data_in(39,50),
			data_out           => s_data_out(39,50),
			out1               => s_out1(39,50),
			out2               => s_out2(39,50),
			lock_lower_row_out => s_locks_lower_out(39,50),
			lock_lower_row_in  => s_locks_lower_in(39,50),
			in1                => s_in1(39,50),
			in2                => s_in2(39,50),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(50)
		);
	s_in1(39,50)            <= s_out1(40,50);
	s_in2(39,50)            <= s_out2(40,51);
	s_locks_lower_in(39,50) <= s_locks_lower_out(40,50);

		normal_cell_39_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,51),
			fetch              => s_fetch(39,51),
			data_in            => s_data_in(39,51),
			data_out           => s_data_out(39,51),
			out1               => s_out1(39,51),
			out2               => s_out2(39,51),
			lock_lower_row_out => s_locks_lower_out(39,51),
			lock_lower_row_in  => s_locks_lower_in(39,51),
			in1                => s_in1(39,51),
			in2                => s_in2(39,51),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(51)
		);
	s_in1(39,51)            <= s_out1(40,51);
	s_in2(39,51)            <= s_out2(40,52);
	s_locks_lower_in(39,51) <= s_locks_lower_out(40,51);

		normal_cell_39_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,52),
			fetch              => s_fetch(39,52),
			data_in            => s_data_in(39,52),
			data_out           => s_data_out(39,52),
			out1               => s_out1(39,52),
			out2               => s_out2(39,52),
			lock_lower_row_out => s_locks_lower_out(39,52),
			lock_lower_row_in  => s_locks_lower_in(39,52),
			in1                => s_in1(39,52),
			in2                => s_in2(39,52),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(52)
		);
	s_in1(39,52)            <= s_out1(40,52);
	s_in2(39,52)            <= s_out2(40,53);
	s_locks_lower_in(39,52) <= s_locks_lower_out(40,52);

		normal_cell_39_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,53),
			fetch              => s_fetch(39,53),
			data_in            => s_data_in(39,53),
			data_out           => s_data_out(39,53),
			out1               => s_out1(39,53),
			out2               => s_out2(39,53),
			lock_lower_row_out => s_locks_lower_out(39,53),
			lock_lower_row_in  => s_locks_lower_in(39,53),
			in1                => s_in1(39,53),
			in2                => s_in2(39,53),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(53)
		);
	s_in1(39,53)            <= s_out1(40,53);
	s_in2(39,53)            <= s_out2(40,54);
	s_locks_lower_in(39,53) <= s_locks_lower_out(40,53);

		normal_cell_39_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,54),
			fetch              => s_fetch(39,54),
			data_in            => s_data_in(39,54),
			data_out           => s_data_out(39,54),
			out1               => s_out1(39,54),
			out2               => s_out2(39,54),
			lock_lower_row_out => s_locks_lower_out(39,54),
			lock_lower_row_in  => s_locks_lower_in(39,54),
			in1                => s_in1(39,54),
			in2                => s_in2(39,54),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(54)
		);
	s_in1(39,54)            <= s_out1(40,54);
	s_in2(39,54)            <= s_out2(40,55);
	s_locks_lower_in(39,54) <= s_locks_lower_out(40,54);

		normal_cell_39_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,55),
			fetch              => s_fetch(39,55),
			data_in            => s_data_in(39,55),
			data_out           => s_data_out(39,55),
			out1               => s_out1(39,55),
			out2               => s_out2(39,55),
			lock_lower_row_out => s_locks_lower_out(39,55),
			lock_lower_row_in  => s_locks_lower_in(39,55),
			in1                => s_in1(39,55),
			in2                => s_in2(39,55),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(55)
		);
	s_in1(39,55)            <= s_out1(40,55);
	s_in2(39,55)            <= s_out2(40,56);
	s_locks_lower_in(39,55) <= s_locks_lower_out(40,55);

		normal_cell_39_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,56),
			fetch              => s_fetch(39,56),
			data_in            => s_data_in(39,56),
			data_out           => s_data_out(39,56),
			out1               => s_out1(39,56),
			out2               => s_out2(39,56),
			lock_lower_row_out => s_locks_lower_out(39,56),
			lock_lower_row_in  => s_locks_lower_in(39,56),
			in1                => s_in1(39,56),
			in2                => s_in2(39,56),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(56)
		);
	s_in1(39,56)            <= s_out1(40,56);
	s_in2(39,56)            <= s_out2(40,57);
	s_locks_lower_in(39,56) <= s_locks_lower_out(40,56);

		normal_cell_39_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,57),
			fetch              => s_fetch(39,57),
			data_in            => s_data_in(39,57),
			data_out           => s_data_out(39,57),
			out1               => s_out1(39,57),
			out2               => s_out2(39,57),
			lock_lower_row_out => s_locks_lower_out(39,57),
			lock_lower_row_in  => s_locks_lower_in(39,57),
			in1                => s_in1(39,57),
			in2                => s_in2(39,57),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(57)
		);
	s_in1(39,57)            <= s_out1(40,57);
	s_in2(39,57)            <= s_out2(40,58);
	s_locks_lower_in(39,57) <= s_locks_lower_out(40,57);

		normal_cell_39_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,58),
			fetch              => s_fetch(39,58),
			data_in            => s_data_in(39,58),
			data_out           => s_data_out(39,58),
			out1               => s_out1(39,58),
			out2               => s_out2(39,58),
			lock_lower_row_out => s_locks_lower_out(39,58),
			lock_lower_row_in  => s_locks_lower_in(39,58),
			in1                => s_in1(39,58),
			in2                => s_in2(39,58),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(58)
		);
	s_in1(39,58)            <= s_out1(40,58);
	s_in2(39,58)            <= s_out2(40,59);
	s_locks_lower_in(39,58) <= s_locks_lower_out(40,58);

		normal_cell_39_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,59),
			fetch              => s_fetch(39,59),
			data_in            => s_data_in(39,59),
			data_out           => s_data_out(39,59),
			out1               => s_out1(39,59),
			out2               => s_out2(39,59),
			lock_lower_row_out => s_locks_lower_out(39,59),
			lock_lower_row_in  => s_locks_lower_in(39,59),
			in1                => s_in1(39,59),
			in2                => s_in2(39,59),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(59)
		);
	s_in1(39,59)            <= s_out1(40,59);
	s_in2(39,59)            <= s_out2(40,60);
	s_locks_lower_in(39,59) <= s_locks_lower_out(40,59);

		last_col_cell_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(39,60),
			fetch              => s_fetch(39,60),
			data_in            => s_data_in(39,60),
			data_out           => s_data_out(39,60),
			out1               => s_out1(39,60),
			out2               => s_out2(39,60),
			lock_lower_row_out => s_locks_lower_out(39,60),
			lock_lower_row_in  => s_locks_lower_in(39,60),
			in1                => s_in1(39,60),
			in2                => (others => '0'),
			lock_row           => s_locks(39),
			piv_found          => s_piv_found,
			row_data           => s_row_data(39),
			col_data           => s_col_data(60)
		);
	s_in1(39,60)            <= s_out1(40,60);
	s_locks_lower_in(39,60) <= s_locks_lower_out(40,60);

		normal_cell_40_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,1),
			fetch              => s_fetch(40,1),
			data_in            => s_data_in(40,1),
			data_out           => s_data_out(40,1),
			out1               => s_out1(40,1),
			out2               => s_out2(40,1),
			lock_lower_row_out => s_locks_lower_out(40,1),
			lock_lower_row_in  => s_locks_lower_in(40,1),
			in1                => s_in1(40,1),
			in2                => s_in2(40,1),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(1)
		);
	s_in1(40,1)            <= s_out1(41,1);
	s_in2(40,1)            <= s_out2(41,2);
	s_locks_lower_in(40,1) <= s_locks_lower_out(41,1);

		normal_cell_40_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,2),
			fetch              => s_fetch(40,2),
			data_in            => s_data_in(40,2),
			data_out           => s_data_out(40,2),
			out1               => s_out1(40,2),
			out2               => s_out2(40,2),
			lock_lower_row_out => s_locks_lower_out(40,2),
			lock_lower_row_in  => s_locks_lower_in(40,2),
			in1                => s_in1(40,2),
			in2                => s_in2(40,2),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(2)
		);
	s_in1(40,2)            <= s_out1(41,2);
	s_in2(40,2)            <= s_out2(41,3);
	s_locks_lower_in(40,2) <= s_locks_lower_out(41,2);

		normal_cell_40_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,3),
			fetch              => s_fetch(40,3),
			data_in            => s_data_in(40,3),
			data_out           => s_data_out(40,3),
			out1               => s_out1(40,3),
			out2               => s_out2(40,3),
			lock_lower_row_out => s_locks_lower_out(40,3),
			lock_lower_row_in  => s_locks_lower_in(40,3),
			in1                => s_in1(40,3),
			in2                => s_in2(40,3),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(3)
		);
	s_in1(40,3)            <= s_out1(41,3);
	s_in2(40,3)            <= s_out2(41,4);
	s_locks_lower_in(40,3) <= s_locks_lower_out(41,3);

		normal_cell_40_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,4),
			fetch              => s_fetch(40,4),
			data_in            => s_data_in(40,4),
			data_out           => s_data_out(40,4),
			out1               => s_out1(40,4),
			out2               => s_out2(40,4),
			lock_lower_row_out => s_locks_lower_out(40,4),
			lock_lower_row_in  => s_locks_lower_in(40,4),
			in1                => s_in1(40,4),
			in2                => s_in2(40,4),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(4)
		);
	s_in1(40,4)            <= s_out1(41,4);
	s_in2(40,4)            <= s_out2(41,5);
	s_locks_lower_in(40,4) <= s_locks_lower_out(41,4);

		normal_cell_40_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,5),
			fetch              => s_fetch(40,5),
			data_in            => s_data_in(40,5),
			data_out           => s_data_out(40,5),
			out1               => s_out1(40,5),
			out2               => s_out2(40,5),
			lock_lower_row_out => s_locks_lower_out(40,5),
			lock_lower_row_in  => s_locks_lower_in(40,5),
			in1                => s_in1(40,5),
			in2                => s_in2(40,5),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(5)
		);
	s_in1(40,5)            <= s_out1(41,5);
	s_in2(40,5)            <= s_out2(41,6);
	s_locks_lower_in(40,5) <= s_locks_lower_out(41,5);

		normal_cell_40_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,6),
			fetch              => s_fetch(40,6),
			data_in            => s_data_in(40,6),
			data_out           => s_data_out(40,6),
			out1               => s_out1(40,6),
			out2               => s_out2(40,6),
			lock_lower_row_out => s_locks_lower_out(40,6),
			lock_lower_row_in  => s_locks_lower_in(40,6),
			in1                => s_in1(40,6),
			in2                => s_in2(40,6),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(6)
		);
	s_in1(40,6)            <= s_out1(41,6);
	s_in2(40,6)            <= s_out2(41,7);
	s_locks_lower_in(40,6) <= s_locks_lower_out(41,6);

		normal_cell_40_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,7),
			fetch              => s_fetch(40,7),
			data_in            => s_data_in(40,7),
			data_out           => s_data_out(40,7),
			out1               => s_out1(40,7),
			out2               => s_out2(40,7),
			lock_lower_row_out => s_locks_lower_out(40,7),
			lock_lower_row_in  => s_locks_lower_in(40,7),
			in1                => s_in1(40,7),
			in2                => s_in2(40,7),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(7)
		);
	s_in1(40,7)            <= s_out1(41,7);
	s_in2(40,7)            <= s_out2(41,8);
	s_locks_lower_in(40,7) <= s_locks_lower_out(41,7);

		normal_cell_40_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,8),
			fetch              => s_fetch(40,8),
			data_in            => s_data_in(40,8),
			data_out           => s_data_out(40,8),
			out1               => s_out1(40,8),
			out2               => s_out2(40,8),
			lock_lower_row_out => s_locks_lower_out(40,8),
			lock_lower_row_in  => s_locks_lower_in(40,8),
			in1                => s_in1(40,8),
			in2                => s_in2(40,8),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(8)
		);
	s_in1(40,8)            <= s_out1(41,8);
	s_in2(40,8)            <= s_out2(41,9);
	s_locks_lower_in(40,8) <= s_locks_lower_out(41,8);

		normal_cell_40_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,9),
			fetch              => s_fetch(40,9),
			data_in            => s_data_in(40,9),
			data_out           => s_data_out(40,9),
			out1               => s_out1(40,9),
			out2               => s_out2(40,9),
			lock_lower_row_out => s_locks_lower_out(40,9),
			lock_lower_row_in  => s_locks_lower_in(40,9),
			in1                => s_in1(40,9),
			in2                => s_in2(40,9),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(9)
		);
	s_in1(40,9)            <= s_out1(41,9);
	s_in2(40,9)            <= s_out2(41,10);
	s_locks_lower_in(40,9) <= s_locks_lower_out(41,9);

		normal_cell_40_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,10),
			fetch              => s_fetch(40,10),
			data_in            => s_data_in(40,10),
			data_out           => s_data_out(40,10),
			out1               => s_out1(40,10),
			out2               => s_out2(40,10),
			lock_lower_row_out => s_locks_lower_out(40,10),
			lock_lower_row_in  => s_locks_lower_in(40,10),
			in1                => s_in1(40,10),
			in2                => s_in2(40,10),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(10)
		);
	s_in1(40,10)            <= s_out1(41,10);
	s_in2(40,10)            <= s_out2(41,11);
	s_locks_lower_in(40,10) <= s_locks_lower_out(41,10);

		normal_cell_40_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,11),
			fetch              => s_fetch(40,11),
			data_in            => s_data_in(40,11),
			data_out           => s_data_out(40,11),
			out1               => s_out1(40,11),
			out2               => s_out2(40,11),
			lock_lower_row_out => s_locks_lower_out(40,11),
			lock_lower_row_in  => s_locks_lower_in(40,11),
			in1                => s_in1(40,11),
			in2                => s_in2(40,11),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(11)
		);
	s_in1(40,11)            <= s_out1(41,11);
	s_in2(40,11)            <= s_out2(41,12);
	s_locks_lower_in(40,11) <= s_locks_lower_out(41,11);

		normal_cell_40_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,12),
			fetch              => s_fetch(40,12),
			data_in            => s_data_in(40,12),
			data_out           => s_data_out(40,12),
			out1               => s_out1(40,12),
			out2               => s_out2(40,12),
			lock_lower_row_out => s_locks_lower_out(40,12),
			lock_lower_row_in  => s_locks_lower_in(40,12),
			in1                => s_in1(40,12),
			in2                => s_in2(40,12),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(12)
		);
	s_in1(40,12)            <= s_out1(41,12);
	s_in2(40,12)            <= s_out2(41,13);
	s_locks_lower_in(40,12) <= s_locks_lower_out(41,12);

		normal_cell_40_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,13),
			fetch              => s_fetch(40,13),
			data_in            => s_data_in(40,13),
			data_out           => s_data_out(40,13),
			out1               => s_out1(40,13),
			out2               => s_out2(40,13),
			lock_lower_row_out => s_locks_lower_out(40,13),
			lock_lower_row_in  => s_locks_lower_in(40,13),
			in1                => s_in1(40,13),
			in2                => s_in2(40,13),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(13)
		);
	s_in1(40,13)            <= s_out1(41,13);
	s_in2(40,13)            <= s_out2(41,14);
	s_locks_lower_in(40,13) <= s_locks_lower_out(41,13);

		normal_cell_40_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,14),
			fetch              => s_fetch(40,14),
			data_in            => s_data_in(40,14),
			data_out           => s_data_out(40,14),
			out1               => s_out1(40,14),
			out2               => s_out2(40,14),
			lock_lower_row_out => s_locks_lower_out(40,14),
			lock_lower_row_in  => s_locks_lower_in(40,14),
			in1                => s_in1(40,14),
			in2                => s_in2(40,14),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(14)
		);
	s_in1(40,14)            <= s_out1(41,14);
	s_in2(40,14)            <= s_out2(41,15);
	s_locks_lower_in(40,14) <= s_locks_lower_out(41,14);

		normal_cell_40_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,15),
			fetch              => s_fetch(40,15),
			data_in            => s_data_in(40,15),
			data_out           => s_data_out(40,15),
			out1               => s_out1(40,15),
			out2               => s_out2(40,15),
			lock_lower_row_out => s_locks_lower_out(40,15),
			lock_lower_row_in  => s_locks_lower_in(40,15),
			in1                => s_in1(40,15),
			in2                => s_in2(40,15),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(15)
		);
	s_in1(40,15)            <= s_out1(41,15);
	s_in2(40,15)            <= s_out2(41,16);
	s_locks_lower_in(40,15) <= s_locks_lower_out(41,15);

		normal_cell_40_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,16),
			fetch              => s_fetch(40,16),
			data_in            => s_data_in(40,16),
			data_out           => s_data_out(40,16),
			out1               => s_out1(40,16),
			out2               => s_out2(40,16),
			lock_lower_row_out => s_locks_lower_out(40,16),
			lock_lower_row_in  => s_locks_lower_in(40,16),
			in1                => s_in1(40,16),
			in2                => s_in2(40,16),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(16)
		);
	s_in1(40,16)            <= s_out1(41,16);
	s_in2(40,16)            <= s_out2(41,17);
	s_locks_lower_in(40,16) <= s_locks_lower_out(41,16);

		normal_cell_40_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,17),
			fetch              => s_fetch(40,17),
			data_in            => s_data_in(40,17),
			data_out           => s_data_out(40,17),
			out1               => s_out1(40,17),
			out2               => s_out2(40,17),
			lock_lower_row_out => s_locks_lower_out(40,17),
			lock_lower_row_in  => s_locks_lower_in(40,17),
			in1                => s_in1(40,17),
			in2                => s_in2(40,17),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(17)
		);
	s_in1(40,17)            <= s_out1(41,17);
	s_in2(40,17)            <= s_out2(41,18);
	s_locks_lower_in(40,17) <= s_locks_lower_out(41,17);

		normal_cell_40_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,18),
			fetch              => s_fetch(40,18),
			data_in            => s_data_in(40,18),
			data_out           => s_data_out(40,18),
			out1               => s_out1(40,18),
			out2               => s_out2(40,18),
			lock_lower_row_out => s_locks_lower_out(40,18),
			lock_lower_row_in  => s_locks_lower_in(40,18),
			in1                => s_in1(40,18),
			in2                => s_in2(40,18),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(18)
		);
	s_in1(40,18)            <= s_out1(41,18);
	s_in2(40,18)            <= s_out2(41,19);
	s_locks_lower_in(40,18) <= s_locks_lower_out(41,18);

		normal_cell_40_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,19),
			fetch              => s_fetch(40,19),
			data_in            => s_data_in(40,19),
			data_out           => s_data_out(40,19),
			out1               => s_out1(40,19),
			out2               => s_out2(40,19),
			lock_lower_row_out => s_locks_lower_out(40,19),
			lock_lower_row_in  => s_locks_lower_in(40,19),
			in1                => s_in1(40,19),
			in2                => s_in2(40,19),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(19)
		);
	s_in1(40,19)            <= s_out1(41,19);
	s_in2(40,19)            <= s_out2(41,20);
	s_locks_lower_in(40,19) <= s_locks_lower_out(41,19);

		normal_cell_40_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,20),
			fetch              => s_fetch(40,20),
			data_in            => s_data_in(40,20),
			data_out           => s_data_out(40,20),
			out1               => s_out1(40,20),
			out2               => s_out2(40,20),
			lock_lower_row_out => s_locks_lower_out(40,20),
			lock_lower_row_in  => s_locks_lower_in(40,20),
			in1                => s_in1(40,20),
			in2                => s_in2(40,20),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(20)
		);
	s_in1(40,20)            <= s_out1(41,20);
	s_in2(40,20)            <= s_out2(41,21);
	s_locks_lower_in(40,20) <= s_locks_lower_out(41,20);

		normal_cell_40_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,21),
			fetch              => s_fetch(40,21),
			data_in            => s_data_in(40,21),
			data_out           => s_data_out(40,21),
			out1               => s_out1(40,21),
			out2               => s_out2(40,21),
			lock_lower_row_out => s_locks_lower_out(40,21),
			lock_lower_row_in  => s_locks_lower_in(40,21),
			in1                => s_in1(40,21),
			in2                => s_in2(40,21),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(21)
		);
	s_in1(40,21)            <= s_out1(41,21);
	s_in2(40,21)            <= s_out2(41,22);
	s_locks_lower_in(40,21) <= s_locks_lower_out(41,21);

		normal_cell_40_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,22),
			fetch              => s_fetch(40,22),
			data_in            => s_data_in(40,22),
			data_out           => s_data_out(40,22),
			out1               => s_out1(40,22),
			out2               => s_out2(40,22),
			lock_lower_row_out => s_locks_lower_out(40,22),
			lock_lower_row_in  => s_locks_lower_in(40,22),
			in1                => s_in1(40,22),
			in2                => s_in2(40,22),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(22)
		);
	s_in1(40,22)            <= s_out1(41,22);
	s_in2(40,22)            <= s_out2(41,23);
	s_locks_lower_in(40,22) <= s_locks_lower_out(41,22);

		normal_cell_40_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,23),
			fetch              => s_fetch(40,23),
			data_in            => s_data_in(40,23),
			data_out           => s_data_out(40,23),
			out1               => s_out1(40,23),
			out2               => s_out2(40,23),
			lock_lower_row_out => s_locks_lower_out(40,23),
			lock_lower_row_in  => s_locks_lower_in(40,23),
			in1                => s_in1(40,23),
			in2                => s_in2(40,23),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(23)
		);
	s_in1(40,23)            <= s_out1(41,23);
	s_in2(40,23)            <= s_out2(41,24);
	s_locks_lower_in(40,23) <= s_locks_lower_out(41,23);

		normal_cell_40_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,24),
			fetch              => s_fetch(40,24),
			data_in            => s_data_in(40,24),
			data_out           => s_data_out(40,24),
			out1               => s_out1(40,24),
			out2               => s_out2(40,24),
			lock_lower_row_out => s_locks_lower_out(40,24),
			lock_lower_row_in  => s_locks_lower_in(40,24),
			in1                => s_in1(40,24),
			in2                => s_in2(40,24),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(24)
		);
	s_in1(40,24)            <= s_out1(41,24);
	s_in2(40,24)            <= s_out2(41,25);
	s_locks_lower_in(40,24) <= s_locks_lower_out(41,24);

		normal_cell_40_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,25),
			fetch              => s_fetch(40,25),
			data_in            => s_data_in(40,25),
			data_out           => s_data_out(40,25),
			out1               => s_out1(40,25),
			out2               => s_out2(40,25),
			lock_lower_row_out => s_locks_lower_out(40,25),
			lock_lower_row_in  => s_locks_lower_in(40,25),
			in1                => s_in1(40,25),
			in2                => s_in2(40,25),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(25)
		);
	s_in1(40,25)            <= s_out1(41,25);
	s_in2(40,25)            <= s_out2(41,26);
	s_locks_lower_in(40,25) <= s_locks_lower_out(41,25);

		normal_cell_40_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,26),
			fetch              => s_fetch(40,26),
			data_in            => s_data_in(40,26),
			data_out           => s_data_out(40,26),
			out1               => s_out1(40,26),
			out2               => s_out2(40,26),
			lock_lower_row_out => s_locks_lower_out(40,26),
			lock_lower_row_in  => s_locks_lower_in(40,26),
			in1                => s_in1(40,26),
			in2                => s_in2(40,26),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(26)
		);
	s_in1(40,26)            <= s_out1(41,26);
	s_in2(40,26)            <= s_out2(41,27);
	s_locks_lower_in(40,26) <= s_locks_lower_out(41,26);

		normal_cell_40_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,27),
			fetch              => s_fetch(40,27),
			data_in            => s_data_in(40,27),
			data_out           => s_data_out(40,27),
			out1               => s_out1(40,27),
			out2               => s_out2(40,27),
			lock_lower_row_out => s_locks_lower_out(40,27),
			lock_lower_row_in  => s_locks_lower_in(40,27),
			in1                => s_in1(40,27),
			in2                => s_in2(40,27),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(27)
		);
	s_in1(40,27)            <= s_out1(41,27);
	s_in2(40,27)            <= s_out2(41,28);
	s_locks_lower_in(40,27) <= s_locks_lower_out(41,27);

		normal_cell_40_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,28),
			fetch              => s_fetch(40,28),
			data_in            => s_data_in(40,28),
			data_out           => s_data_out(40,28),
			out1               => s_out1(40,28),
			out2               => s_out2(40,28),
			lock_lower_row_out => s_locks_lower_out(40,28),
			lock_lower_row_in  => s_locks_lower_in(40,28),
			in1                => s_in1(40,28),
			in2                => s_in2(40,28),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(28)
		);
	s_in1(40,28)            <= s_out1(41,28);
	s_in2(40,28)            <= s_out2(41,29);
	s_locks_lower_in(40,28) <= s_locks_lower_out(41,28);

		normal_cell_40_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,29),
			fetch              => s_fetch(40,29),
			data_in            => s_data_in(40,29),
			data_out           => s_data_out(40,29),
			out1               => s_out1(40,29),
			out2               => s_out2(40,29),
			lock_lower_row_out => s_locks_lower_out(40,29),
			lock_lower_row_in  => s_locks_lower_in(40,29),
			in1                => s_in1(40,29),
			in2                => s_in2(40,29),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(29)
		);
	s_in1(40,29)            <= s_out1(41,29);
	s_in2(40,29)            <= s_out2(41,30);
	s_locks_lower_in(40,29) <= s_locks_lower_out(41,29);

		normal_cell_40_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,30),
			fetch              => s_fetch(40,30),
			data_in            => s_data_in(40,30),
			data_out           => s_data_out(40,30),
			out1               => s_out1(40,30),
			out2               => s_out2(40,30),
			lock_lower_row_out => s_locks_lower_out(40,30),
			lock_lower_row_in  => s_locks_lower_in(40,30),
			in1                => s_in1(40,30),
			in2                => s_in2(40,30),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(30)
		);
	s_in1(40,30)            <= s_out1(41,30);
	s_in2(40,30)            <= s_out2(41,31);
	s_locks_lower_in(40,30) <= s_locks_lower_out(41,30);

		normal_cell_40_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,31),
			fetch              => s_fetch(40,31),
			data_in            => s_data_in(40,31),
			data_out           => s_data_out(40,31),
			out1               => s_out1(40,31),
			out2               => s_out2(40,31),
			lock_lower_row_out => s_locks_lower_out(40,31),
			lock_lower_row_in  => s_locks_lower_in(40,31),
			in1                => s_in1(40,31),
			in2                => s_in2(40,31),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(31)
		);
	s_in1(40,31)            <= s_out1(41,31);
	s_in2(40,31)            <= s_out2(41,32);
	s_locks_lower_in(40,31) <= s_locks_lower_out(41,31);

		normal_cell_40_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,32),
			fetch              => s_fetch(40,32),
			data_in            => s_data_in(40,32),
			data_out           => s_data_out(40,32),
			out1               => s_out1(40,32),
			out2               => s_out2(40,32),
			lock_lower_row_out => s_locks_lower_out(40,32),
			lock_lower_row_in  => s_locks_lower_in(40,32),
			in1                => s_in1(40,32),
			in2                => s_in2(40,32),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(32)
		);
	s_in1(40,32)            <= s_out1(41,32);
	s_in2(40,32)            <= s_out2(41,33);
	s_locks_lower_in(40,32) <= s_locks_lower_out(41,32);

		normal_cell_40_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,33),
			fetch              => s_fetch(40,33),
			data_in            => s_data_in(40,33),
			data_out           => s_data_out(40,33),
			out1               => s_out1(40,33),
			out2               => s_out2(40,33),
			lock_lower_row_out => s_locks_lower_out(40,33),
			lock_lower_row_in  => s_locks_lower_in(40,33),
			in1                => s_in1(40,33),
			in2                => s_in2(40,33),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(33)
		);
	s_in1(40,33)            <= s_out1(41,33);
	s_in2(40,33)            <= s_out2(41,34);
	s_locks_lower_in(40,33) <= s_locks_lower_out(41,33);

		normal_cell_40_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,34),
			fetch              => s_fetch(40,34),
			data_in            => s_data_in(40,34),
			data_out           => s_data_out(40,34),
			out1               => s_out1(40,34),
			out2               => s_out2(40,34),
			lock_lower_row_out => s_locks_lower_out(40,34),
			lock_lower_row_in  => s_locks_lower_in(40,34),
			in1                => s_in1(40,34),
			in2                => s_in2(40,34),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(34)
		);
	s_in1(40,34)            <= s_out1(41,34);
	s_in2(40,34)            <= s_out2(41,35);
	s_locks_lower_in(40,34) <= s_locks_lower_out(41,34);

		normal_cell_40_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,35),
			fetch              => s_fetch(40,35),
			data_in            => s_data_in(40,35),
			data_out           => s_data_out(40,35),
			out1               => s_out1(40,35),
			out2               => s_out2(40,35),
			lock_lower_row_out => s_locks_lower_out(40,35),
			lock_lower_row_in  => s_locks_lower_in(40,35),
			in1                => s_in1(40,35),
			in2                => s_in2(40,35),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(35)
		);
	s_in1(40,35)            <= s_out1(41,35);
	s_in2(40,35)            <= s_out2(41,36);
	s_locks_lower_in(40,35) <= s_locks_lower_out(41,35);

		normal_cell_40_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,36),
			fetch              => s_fetch(40,36),
			data_in            => s_data_in(40,36),
			data_out           => s_data_out(40,36),
			out1               => s_out1(40,36),
			out2               => s_out2(40,36),
			lock_lower_row_out => s_locks_lower_out(40,36),
			lock_lower_row_in  => s_locks_lower_in(40,36),
			in1                => s_in1(40,36),
			in2                => s_in2(40,36),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(36)
		);
	s_in1(40,36)            <= s_out1(41,36);
	s_in2(40,36)            <= s_out2(41,37);
	s_locks_lower_in(40,36) <= s_locks_lower_out(41,36);

		normal_cell_40_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,37),
			fetch              => s_fetch(40,37),
			data_in            => s_data_in(40,37),
			data_out           => s_data_out(40,37),
			out1               => s_out1(40,37),
			out2               => s_out2(40,37),
			lock_lower_row_out => s_locks_lower_out(40,37),
			lock_lower_row_in  => s_locks_lower_in(40,37),
			in1                => s_in1(40,37),
			in2                => s_in2(40,37),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(37)
		);
	s_in1(40,37)            <= s_out1(41,37);
	s_in2(40,37)            <= s_out2(41,38);
	s_locks_lower_in(40,37) <= s_locks_lower_out(41,37);

		normal_cell_40_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,38),
			fetch              => s_fetch(40,38),
			data_in            => s_data_in(40,38),
			data_out           => s_data_out(40,38),
			out1               => s_out1(40,38),
			out2               => s_out2(40,38),
			lock_lower_row_out => s_locks_lower_out(40,38),
			lock_lower_row_in  => s_locks_lower_in(40,38),
			in1                => s_in1(40,38),
			in2                => s_in2(40,38),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(38)
		);
	s_in1(40,38)            <= s_out1(41,38);
	s_in2(40,38)            <= s_out2(41,39);
	s_locks_lower_in(40,38) <= s_locks_lower_out(41,38);

		normal_cell_40_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,39),
			fetch              => s_fetch(40,39),
			data_in            => s_data_in(40,39),
			data_out           => s_data_out(40,39),
			out1               => s_out1(40,39),
			out2               => s_out2(40,39),
			lock_lower_row_out => s_locks_lower_out(40,39),
			lock_lower_row_in  => s_locks_lower_in(40,39),
			in1                => s_in1(40,39),
			in2                => s_in2(40,39),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(39)
		);
	s_in1(40,39)            <= s_out1(41,39);
	s_in2(40,39)            <= s_out2(41,40);
	s_locks_lower_in(40,39) <= s_locks_lower_out(41,39);

		normal_cell_40_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,40),
			fetch              => s_fetch(40,40),
			data_in            => s_data_in(40,40),
			data_out           => s_data_out(40,40),
			out1               => s_out1(40,40),
			out2               => s_out2(40,40),
			lock_lower_row_out => s_locks_lower_out(40,40),
			lock_lower_row_in  => s_locks_lower_in(40,40),
			in1                => s_in1(40,40),
			in2                => s_in2(40,40),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(40)
		);
	s_in1(40,40)            <= s_out1(41,40);
	s_in2(40,40)            <= s_out2(41,41);
	s_locks_lower_in(40,40) <= s_locks_lower_out(41,40);

		normal_cell_40_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,41),
			fetch              => s_fetch(40,41),
			data_in            => s_data_in(40,41),
			data_out           => s_data_out(40,41),
			out1               => s_out1(40,41),
			out2               => s_out2(40,41),
			lock_lower_row_out => s_locks_lower_out(40,41),
			lock_lower_row_in  => s_locks_lower_in(40,41),
			in1                => s_in1(40,41),
			in2                => s_in2(40,41),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(41)
		);
	s_in1(40,41)            <= s_out1(41,41);
	s_in2(40,41)            <= s_out2(41,42);
	s_locks_lower_in(40,41) <= s_locks_lower_out(41,41);

		normal_cell_40_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,42),
			fetch              => s_fetch(40,42),
			data_in            => s_data_in(40,42),
			data_out           => s_data_out(40,42),
			out1               => s_out1(40,42),
			out2               => s_out2(40,42),
			lock_lower_row_out => s_locks_lower_out(40,42),
			lock_lower_row_in  => s_locks_lower_in(40,42),
			in1                => s_in1(40,42),
			in2                => s_in2(40,42),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(42)
		);
	s_in1(40,42)            <= s_out1(41,42);
	s_in2(40,42)            <= s_out2(41,43);
	s_locks_lower_in(40,42) <= s_locks_lower_out(41,42);

		normal_cell_40_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,43),
			fetch              => s_fetch(40,43),
			data_in            => s_data_in(40,43),
			data_out           => s_data_out(40,43),
			out1               => s_out1(40,43),
			out2               => s_out2(40,43),
			lock_lower_row_out => s_locks_lower_out(40,43),
			lock_lower_row_in  => s_locks_lower_in(40,43),
			in1                => s_in1(40,43),
			in2                => s_in2(40,43),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(43)
		);
	s_in1(40,43)            <= s_out1(41,43);
	s_in2(40,43)            <= s_out2(41,44);
	s_locks_lower_in(40,43) <= s_locks_lower_out(41,43);

		normal_cell_40_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,44),
			fetch              => s_fetch(40,44),
			data_in            => s_data_in(40,44),
			data_out           => s_data_out(40,44),
			out1               => s_out1(40,44),
			out2               => s_out2(40,44),
			lock_lower_row_out => s_locks_lower_out(40,44),
			lock_lower_row_in  => s_locks_lower_in(40,44),
			in1                => s_in1(40,44),
			in2                => s_in2(40,44),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(44)
		);
	s_in1(40,44)            <= s_out1(41,44);
	s_in2(40,44)            <= s_out2(41,45);
	s_locks_lower_in(40,44) <= s_locks_lower_out(41,44);

		normal_cell_40_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,45),
			fetch              => s_fetch(40,45),
			data_in            => s_data_in(40,45),
			data_out           => s_data_out(40,45),
			out1               => s_out1(40,45),
			out2               => s_out2(40,45),
			lock_lower_row_out => s_locks_lower_out(40,45),
			lock_lower_row_in  => s_locks_lower_in(40,45),
			in1                => s_in1(40,45),
			in2                => s_in2(40,45),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(45)
		);
	s_in1(40,45)            <= s_out1(41,45);
	s_in2(40,45)            <= s_out2(41,46);
	s_locks_lower_in(40,45) <= s_locks_lower_out(41,45);

		normal_cell_40_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,46),
			fetch              => s_fetch(40,46),
			data_in            => s_data_in(40,46),
			data_out           => s_data_out(40,46),
			out1               => s_out1(40,46),
			out2               => s_out2(40,46),
			lock_lower_row_out => s_locks_lower_out(40,46),
			lock_lower_row_in  => s_locks_lower_in(40,46),
			in1                => s_in1(40,46),
			in2                => s_in2(40,46),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(46)
		);
	s_in1(40,46)            <= s_out1(41,46);
	s_in2(40,46)            <= s_out2(41,47);
	s_locks_lower_in(40,46) <= s_locks_lower_out(41,46);

		normal_cell_40_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,47),
			fetch              => s_fetch(40,47),
			data_in            => s_data_in(40,47),
			data_out           => s_data_out(40,47),
			out1               => s_out1(40,47),
			out2               => s_out2(40,47),
			lock_lower_row_out => s_locks_lower_out(40,47),
			lock_lower_row_in  => s_locks_lower_in(40,47),
			in1                => s_in1(40,47),
			in2                => s_in2(40,47),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(47)
		);
	s_in1(40,47)            <= s_out1(41,47);
	s_in2(40,47)            <= s_out2(41,48);
	s_locks_lower_in(40,47) <= s_locks_lower_out(41,47);

		normal_cell_40_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,48),
			fetch              => s_fetch(40,48),
			data_in            => s_data_in(40,48),
			data_out           => s_data_out(40,48),
			out1               => s_out1(40,48),
			out2               => s_out2(40,48),
			lock_lower_row_out => s_locks_lower_out(40,48),
			lock_lower_row_in  => s_locks_lower_in(40,48),
			in1                => s_in1(40,48),
			in2                => s_in2(40,48),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(48)
		);
	s_in1(40,48)            <= s_out1(41,48);
	s_in2(40,48)            <= s_out2(41,49);
	s_locks_lower_in(40,48) <= s_locks_lower_out(41,48);

		normal_cell_40_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,49),
			fetch              => s_fetch(40,49),
			data_in            => s_data_in(40,49),
			data_out           => s_data_out(40,49),
			out1               => s_out1(40,49),
			out2               => s_out2(40,49),
			lock_lower_row_out => s_locks_lower_out(40,49),
			lock_lower_row_in  => s_locks_lower_in(40,49),
			in1                => s_in1(40,49),
			in2                => s_in2(40,49),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(49)
		);
	s_in1(40,49)            <= s_out1(41,49);
	s_in2(40,49)            <= s_out2(41,50);
	s_locks_lower_in(40,49) <= s_locks_lower_out(41,49);

		normal_cell_40_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,50),
			fetch              => s_fetch(40,50),
			data_in            => s_data_in(40,50),
			data_out           => s_data_out(40,50),
			out1               => s_out1(40,50),
			out2               => s_out2(40,50),
			lock_lower_row_out => s_locks_lower_out(40,50),
			lock_lower_row_in  => s_locks_lower_in(40,50),
			in1                => s_in1(40,50),
			in2                => s_in2(40,50),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(50)
		);
	s_in1(40,50)            <= s_out1(41,50);
	s_in2(40,50)            <= s_out2(41,51);
	s_locks_lower_in(40,50) <= s_locks_lower_out(41,50);

		normal_cell_40_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,51),
			fetch              => s_fetch(40,51),
			data_in            => s_data_in(40,51),
			data_out           => s_data_out(40,51),
			out1               => s_out1(40,51),
			out2               => s_out2(40,51),
			lock_lower_row_out => s_locks_lower_out(40,51),
			lock_lower_row_in  => s_locks_lower_in(40,51),
			in1                => s_in1(40,51),
			in2                => s_in2(40,51),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(51)
		);
	s_in1(40,51)            <= s_out1(41,51);
	s_in2(40,51)            <= s_out2(41,52);
	s_locks_lower_in(40,51) <= s_locks_lower_out(41,51);

		normal_cell_40_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,52),
			fetch              => s_fetch(40,52),
			data_in            => s_data_in(40,52),
			data_out           => s_data_out(40,52),
			out1               => s_out1(40,52),
			out2               => s_out2(40,52),
			lock_lower_row_out => s_locks_lower_out(40,52),
			lock_lower_row_in  => s_locks_lower_in(40,52),
			in1                => s_in1(40,52),
			in2                => s_in2(40,52),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(52)
		);
	s_in1(40,52)            <= s_out1(41,52);
	s_in2(40,52)            <= s_out2(41,53);
	s_locks_lower_in(40,52) <= s_locks_lower_out(41,52);

		normal_cell_40_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,53),
			fetch              => s_fetch(40,53),
			data_in            => s_data_in(40,53),
			data_out           => s_data_out(40,53),
			out1               => s_out1(40,53),
			out2               => s_out2(40,53),
			lock_lower_row_out => s_locks_lower_out(40,53),
			lock_lower_row_in  => s_locks_lower_in(40,53),
			in1                => s_in1(40,53),
			in2                => s_in2(40,53),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(53)
		);
	s_in1(40,53)            <= s_out1(41,53);
	s_in2(40,53)            <= s_out2(41,54);
	s_locks_lower_in(40,53) <= s_locks_lower_out(41,53);

		normal_cell_40_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,54),
			fetch              => s_fetch(40,54),
			data_in            => s_data_in(40,54),
			data_out           => s_data_out(40,54),
			out1               => s_out1(40,54),
			out2               => s_out2(40,54),
			lock_lower_row_out => s_locks_lower_out(40,54),
			lock_lower_row_in  => s_locks_lower_in(40,54),
			in1                => s_in1(40,54),
			in2                => s_in2(40,54),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(54)
		);
	s_in1(40,54)            <= s_out1(41,54);
	s_in2(40,54)            <= s_out2(41,55);
	s_locks_lower_in(40,54) <= s_locks_lower_out(41,54);

		normal_cell_40_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,55),
			fetch              => s_fetch(40,55),
			data_in            => s_data_in(40,55),
			data_out           => s_data_out(40,55),
			out1               => s_out1(40,55),
			out2               => s_out2(40,55),
			lock_lower_row_out => s_locks_lower_out(40,55),
			lock_lower_row_in  => s_locks_lower_in(40,55),
			in1                => s_in1(40,55),
			in2                => s_in2(40,55),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(55)
		);
	s_in1(40,55)            <= s_out1(41,55);
	s_in2(40,55)            <= s_out2(41,56);
	s_locks_lower_in(40,55) <= s_locks_lower_out(41,55);

		normal_cell_40_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,56),
			fetch              => s_fetch(40,56),
			data_in            => s_data_in(40,56),
			data_out           => s_data_out(40,56),
			out1               => s_out1(40,56),
			out2               => s_out2(40,56),
			lock_lower_row_out => s_locks_lower_out(40,56),
			lock_lower_row_in  => s_locks_lower_in(40,56),
			in1                => s_in1(40,56),
			in2                => s_in2(40,56),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(56)
		);
	s_in1(40,56)            <= s_out1(41,56);
	s_in2(40,56)            <= s_out2(41,57);
	s_locks_lower_in(40,56) <= s_locks_lower_out(41,56);

		normal_cell_40_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,57),
			fetch              => s_fetch(40,57),
			data_in            => s_data_in(40,57),
			data_out           => s_data_out(40,57),
			out1               => s_out1(40,57),
			out2               => s_out2(40,57),
			lock_lower_row_out => s_locks_lower_out(40,57),
			lock_lower_row_in  => s_locks_lower_in(40,57),
			in1                => s_in1(40,57),
			in2                => s_in2(40,57),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(57)
		);
	s_in1(40,57)            <= s_out1(41,57);
	s_in2(40,57)            <= s_out2(41,58);
	s_locks_lower_in(40,57) <= s_locks_lower_out(41,57);

		normal_cell_40_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,58),
			fetch              => s_fetch(40,58),
			data_in            => s_data_in(40,58),
			data_out           => s_data_out(40,58),
			out1               => s_out1(40,58),
			out2               => s_out2(40,58),
			lock_lower_row_out => s_locks_lower_out(40,58),
			lock_lower_row_in  => s_locks_lower_in(40,58),
			in1                => s_in1(40,58),
			in2                => s_in2(40,58),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(58)
		);
	s_in1(40,58)            <= s_out1(41,58);
	s_in2(40,58)            <= s_out2(41,59);
	s_locks_lower_in(40,58) <= s_locks_lower_out(41,58);

		normal_cell_40_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,59),
			fetch              => s_fetch(40,59),
			data_in            => s_data_in(40,59),
			data_out           => s_data_out(40,59),
			out1               => s_out1(40,59),
			out2               => s_out2(40,59),
			lock_lower_row_out => s_locks_lower_out(40,59),
			lock_lower_row_in  => s_locks_lower_in(40,59),
			in1                => s_in1(40,59),
			in2                => s_in2(40,59),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(59)
		);
	s_in1(40,59)            <= s_out1(41,59);
	s_in2(40,59)            <= s_out2(41,60);
	s_locks_lower_in(40,59) <= s_locks_lower_out(41,59);

		last_col_cell_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(40,60),
			fetch              => s_fetch(40,60),
			data_in            => s_data_in(40,60),
			data_out           => s_data_out(40,60),
			out1               => s_out1(40,60),
			out2               => s_out2(40,60),
			lock_lower_row_out => s_locks_lower_out(40,60),
			lock_lower_row_in  => s_locks_lower_in(40,60),
			in1                => s_in1(40,60),
			in2                => (others => '0'),
			lock_row           => s_locks(40),
			piv_found          => s_piv_found,
			row_data           => s_row_data(40),
			col_data           => s_col_data(60)
		);
	s_in1(40,60)            <= s_out1(41,60);
	s_locks_lower_in(40,60) <= s_locks_lower_out(41,60);

		normal_cell_41_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,1),
			fetch              => s_fetch(41,1),
			data_in            => s_data_in(41,1),
			data_out           => s_data_out(41,1),
			out1               => s_out1(41,1),
			out2               => s_out2(41,1),
			lock_lower_row_out => s_locks_lower_out(41,1),
			lock_lower_row_in  => s_locks_lower_in(41,1),
			in1                => s_in1(41,1),
			in2                => s_in2(41,1),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(1)
		);
	s_in1(41,1)            <= s_out1(42,1);
	s_in2(41,1)            <= s_out2(42,2);
	s_locks_lower_in(41,1) <= s_locks_lower_out(42,1);

		normal_cell_41_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,2),
			fetch              => s_fetch(41,2),
			data_in            => s_data_in(41,2),
			data_out           => s_data_out(41,2),
			out1               => s_out1(41,2),
			out2               => s_out2(41,2),
			lock_lower_row_out => s_locks_lower_out(41,2),
			lock_lower_row_in  => s_locks_lower_in(41,2),
			in1                => s_in1(41,2),
			in2                => s_in2(41,2),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(2)
		);
	s_in1(41,2)            <= s_out1(42,2);
	s_in2(41,2)            <= s_out2(42,3);
	s_locks_lower_in(41,2) <= s_locks_lower_out(42,2);

		normal_cell_41_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,3),
			fetch              => s_fetch(41,3),
			data_in            => s_data_in(41,3),
			data_out           => s_data_out(41,3),
			out1               => s_out1(41,3),
			out2               => s_out2(41,3),
			lock_lower_row_out => s_locks_lower_out(41,3),
			lock_lower_row_in  => s_locks_lower_in(41,3),
			in1                => s_in1(41,3),
			in2                => s_in2(41,3),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(3)
		);
	s_in1(41,3)            <= s_out1(42,3);
	s_in2(41,3)            <= s_out2(42,4);
	s_locks_lower_in(41,3) <= s_locks_lower_out(42,3);

		normal_cell_41_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,4),
			fetch              => s_fetch(41,4),
			data_in            => s_data_in(41,4),
			data_out           => s_data_out(41,4),
			out1               => s_out1(41,4),
			out2               => s_out2(41,4),
			lock_lower_row_out => s_locks_lower_out(41,4),
			lock_lower_row_in  => s_locks_lower_in(41,4),
			in1                => s_in1(41,4),
			in2                => s_in2(41,4),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(4)
		);
	s_in1(41,4)            <= s_out1(42,4);
	s_in2(41,4)            <= s_out2(42,5);
	s_locks_lower_in(41,4) <= s_locks_lower_out(42,4);

		normal_cell_41_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,5),
			fetch              => s_fetch(41,5),
			data_in            => s_data_in(41,5),
			data_out           => s_data_out(41,5),
			out1               => s_out1(41,5),
			out2               => s_out2(41,5),
			lock_lower_row_out => s_locks_lower_out(41,5),
			lock_lower_row_in  => s_locks_lower_in(41,5),
			in1                => s_in1(41,5),
			in2                => s_in2(41,5),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(5)
		);
	s_in1(41,5)            <= s_out1(42,5);
	s_in2(41,5)            <= s_out2(42,6);
	s_locks_lower_in(41,5) <= s_locks_lower_out(42,5);

		normal_cell_41_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,6),
			fetch              => s_fetch(41,6),
			data_in            => s_data_in(41,6),
			data_out           => s_data_out(41,6),
			out1               => s_out1(41,6),
			out2               => s_out2(41,6),
			lock_lower_row_out => s_locks_lower_out(41,6),
			lock_lower_row_in  => s_locks_lower_in(41,6),
			in1                => s_in1(41,6),
			in2                => s_in2(41,6),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(6)
		);
	s_in1(41,6)            <= s_out1(42,6);
	s_in2(41,6)            <= s_out2(42,7);
	s_locks_lower_in(41,6) <= s_locks_lower_out(42,6);

		normal_cell_41_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,7),
			fetch              => s_fetch(41,7),
			data_in            => s_data_in(41,7),
			data_out           => s_data_out(41,7),
			out1               => s_out1(41,7),
			out2               => s_out2(41,7),
			lock_lower_row_out => s_locks_lower_out(41,7),
			lock_lower_row_in  => s_locks_lower_in(41,7),
			in1                => s_in1(41,7),
			in2                => s_in2(41,7),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(7)
		);
	s_in1(41,7)            <= s_out1(42,7);
	s_in2(41,7)            <= s_out2(42,8);
	s_locks_lower_in(41,7) <= s_locks_lower_out(42,7);

		normal_cell_41_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,8),
			fetch              => s_fetch(41,8),
			data_in            => s_data_in(41,8),
			data_out           => s_data_out(41,8),
			out1               => s_out1(41,8),
			out2               => s_out2(41,8),
			lock_lower_row_out => s_locks_lower_out(41,8),
			lock_lower_row_in  => s_locks_lower_in(41,8),
			in1                => s_in1(41,8),
			in2                => s_in2(41,8),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(8)
		);
	s_in1(41,8)            <= s_out1(42,8);
	s_in2(41,8)            <= s_out2(42,9);
	s_locks_lower_in(41,8) <= s_locks_lower_out(42,8);

		normal_cell_41_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,9),
			fetch              => s_fetch(41,9),
			data_in            => s_data_in(41,9),
			data_out           => s_data_out(41,9),
			out1               => s_out1(41,9),
			out2               => s_out2(41,9),
			lock_lower_row_out => s_locks_lower_out(41,9),
			lock_lower_row_in  => s_locks_lower_in(41,9),
			in1                => s_in1(41,9),
			in2                => s_in2(41,9),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(9)
		);
	s_in1(41,9)            <= s_out1(42,9);
	s_in2(41,9)            <= s_out2(42,10);
	s_locks_lower_in(41,9) <= s_locks_lower_out(42,9);

		normal_cell_41_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,10),
			fetch              => s_fetch(41,10),
			data_in            => s_data_in(41,10),
			data_out           => s_data_out(41,10),
			out1               => s_out1(41,10),
			out2               => s_out2(41,10),
			lock_lower_row_out => s_locks_lower_out(41,10),
			lock_lower_row_in  => s_locks_lower_in(41,10),
			in1                => s_in1(41,10),
			in2                => s_in2(41,10),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(10)
		);
	s_in1(41,10)            <= s_out1(42,10);
	s_in2(41,10)            <= s_out2(42,11);
	s_locks_lower_in(41,10) <= s_locks_lower_out(42,10);

		normal_cell_41_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,11),
			fetch              => s_fetch(41,11),
			data_in            => s_data_in(41,11),
			data_out           => s_data_out(41,11),
			out1               => s_out1(41,11),
			out2               => s_out2(41,11),
			lock_lower_row_out => s_locks_lower_out(41,11),
			lock_lower_row_in  => s_locks_lower_in(41,11),
			in1                => s_in1(41,11),
			in2                => s_in2(41,11),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(11)
		);
	s_in1(41,11)            <= s_out1(42,11);
	s_in2(41,11)            <= s_out2(42,12);
	s_locks_lower_in(41,11) <= s_locks_lower_out(42,11);

		normal_cell_41_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,12),
			fetch              => s_fetch(41,12),
			data_in            => s_data_in(41,12),
			data_out           => s_data_out(41,12),
			out1               => s_out1(41,12),
			out2               => s_out2(41,12),
			lock_lower_row_out => s_locks_lower_out(41,12),
			lock_lower_row_in  => s_locks_lower_in(41,12),
			in1                => s_in1(41,12),
			in2                => s_in2(41,12),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(12)
		);
	s_in1(41,12)            <= s_out1(42,12);
	s_in2(41,12)            <= s_out2(42,13);
	s_locks_lower_in(41,12) <= s_locks_lower_out(42,12);

		normal_cell_41_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,13),
			fetch              => s_fetch(41,13),
			data_in            => s_data_in(41,13),
			data_out           => s_data_out(41,13),
			out1               => s_out1(41,13),
			out2               => s_out2(41,13),
			lock_lower_row_out => s_locks_lower_out(41,13),
			lock_lower_row_in  => s_locks_lower_in(41,13),
			in1                => s_in1(41,13),
			in2                => s_in2(41,13),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(13)
		);
	s_in1(41,13)            <= s_out1(42,13);
	s_in2(41,13)            <= s_out2(42,14);
	s_locks_lower_in(41,13) <= s_locks_lower_out(42,13);

		normal_cell_41_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,14),
			fetch              => s_fetch(41,14),
			data_in            => s_data_in(41,14),
			data_out           => s_data_out(41,14),
			out1               => s_out1(41,14),
			out2               => s_out2(41,14),
			lock_lower_row_out => s_locks_lower_out(41,14),
			lock_lower_row_in  => s_locks_lower_in(41,14),
			in1                => s_in1(41,14),
			in2                => s_in2(41,14),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(14)
		);
	s_in1(41,14)            <= s_out1(42,14);
	s_in2(41,14)            <= s_out2(42,15);
	s_locks_lower_in(41,14) <= s_locks_lower_out(42,14);

		normal_cell_41_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,15),
			fetch              => s_fetch(41,15),
			data_in            => s_data_in(41,15),
			data_out           => s_data_out(41,15),
			out1               => s_out1(41,15),
			out2               => s_out2(41,15),
			lock_lower_row_out => s_locks_lower_out(41,15),
			lock_lower_row_in  => s_locks_lower_in(41,15),
			in1                => s_in1(41,15),
			in2                => s_in2(41,15),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(15)
		);
	s_in1(41,15)            <= s_out1(42,15);
	s_in2(41,15)            <= s_out2(42,16);
	s_locks_lower_in(41,15) <= s_locks_lower_out(42,15);

		normal_cell_41_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,16),
			fetch              => s_fetch(41,16),
			data_in            => s_data_in(41,16),
			data_out           => s_data_out(41,16),
			out1               => s_out1(41,16),
			out2               => s_out2(41,16),
			lock_lower_row_out => s_locks_lower_out(41,16),
			lock_lower_row_in  => s_locks_lower_in(41,16),
			in1                => s_in1(41,16),
			in2                => s_in2(41,16),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(16)
		);
	s_in1(41,16)            <= s_out1(42,16);
	s_in2(41,16)            <= s_out2(42,17);
	s_locks_lower_in(41,16) <= s_locks_lower_out(42,16);

		normal_cell_41_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,17),
			fetch              => s_fetch(41,17),
			data_in            => s_data_in(41,17),
			data_out           => s_data_out(41,17),
			out1               => s_out1(41,17),
			out2               => s_out2(41,17),
			lock_lower_row_out => s_locks_lower_out(41,17),
			lock_lower_row_in  => s_locks_lower_in(41,17),
			in1                => s_in1(41,17),
			in2                => s_in2(41,17),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(17)
		);
	s_in1(41,17)            <= s_out1(42,17);
	s_in2(41,17)            <= s_out2(42,18);
	s_locks_lower_in(41,17) <= s_locks_lower_out(42,17);

		normal_cell_41_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,18),
			fetch              => s_fetch(41,18),
			data_in            => s_data_in(41,18),
			data_out           => s_data_out(41,18),
			out1               => s_out1(41,18),
			out2               => s_out2(41,18),
			lock_lower_row_out => s_locks_lower_out(41,18),
			lock_lower_row_in  => s_locks_lower_in(41,18),
			in1                => s_in1(41,18),
			in2                => s_in2(41,18),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(18)
		);
	s_in1(41,18)            <= s_out1(42,18);
	s_in2(41,18)            <= s_out2(42,19);
	s_locks_lower_in(41,18) <= s_locks_lower_out(42,18);

		normal_cell_41_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,19),
			fetch              => s_fetch(41,19),
			data_in            => s_data_in(41,19),
			data_out           => s_data_out(41,19),
			out1               => s_out1(41,19),
			out2               => s_out2(41,19),
			lock_lower_row_out => s_locks_lower_out(41,19),
			lock_lower_row_in  => s_locks_lower_in(41,19),
			in1                => s_in1(41,19),
			in2                => s_in2(41,19),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(19)
		);
	s_in1(41,19)            <= s_out1(42,19);
	s_in2(41,19)            <= s_out2(42,20);
	s_locks_lower_in(41,19) <= s_locks_lower_out(42,19);

		normal_cell_41_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,20),
			fetch              => s_fetch(41,20),
			data_in            => s_data_in(41,20),
			data_out           => s_data_out(41,20),
			out1               => s_out1(41,20),
			out2               => s_out2(41,20),
			lock_lower_row_out => s_locks_lower_out(41,20),
			lock_lower_row_in  => s_locks_lower_in(41,20),
			in1                => s_in1(41,20),
			in2                => s_in2(41,20),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(20)
		);
	s_in1(41,20)            <= s_out1(42,20);
	s_in2(41,20)            <= s_out2(42,21);
	s_locks_lower_in(41,20) <= s_locks_lower_out(42,20);

		normal_cell_41_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,21),
			fetch              => s_fetch(41,21),
			data_in            => s_data_in(41,21),
			data_out           => s_data_out(41,21),
			out1               => s_out1(41,21),
			out2               => s_out2(41,21),
			lock_lower_row_out => s_locks_lower_out(41,21),
			lock_lower_row_in  => s_locks_lower_in(41,21),
			in1                => s_in1(41,21),
			in2                => s_in2(41,21),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(21)
		);
	s_in1(41,21)            <= s_out1(42,21);
	s_in2(41,21)            <= s_out2(42,22);
	s_locks_lower_in(41,21) <= s_locks_lower_out(42,21);

		normal_cell_41_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,22),
			fetch              => s_fetch(41,22),
			data_in            => s_data_in(41,22),
			data_out           => s_data_out(41,22),
			out1               => s_out1(41,22),
			out2               => s_out2(41,22),
			lock_lower_row_out => s_locks_lower_out(41,22),
			lock_lower_row_in  => s_locks_lower_in(41,22),
			in1                => s_in1(41,22),
			in2                => s_in2(41,22),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(22)
		);
	s_in1(41,22)            <= s_out1(42,22);
	s_in2(41,22)            <= s_out2(42,23);
	s_locks_lower_in(41,22) <= s_locks_lower_out(42,22);

		normal_cell_41_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,23),
			fetch              => s_fetch(41,23),
			data_in            => s_data_in(41,23),
			data_out           => s_data_out(41,23),
			out1               => s_out1(41,23),
			out2               => s_out2(41,23),
			lock_lower_row_out => s_locks_lower_out(41,23),
			lock_lower_row_in  => s_locks_lower_in(41,23),
			in1                => s_in1(41,23),
			in2                => s_in2(41,23),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(23)
		);
	s_in1(41,23)            <= s_out1(42,23);
	s_in2(41,23)            <= s_out2(42,24);
	s_locks_lower_in(41,23) <= s_locks_lower_out(42,23);

		normal_cell_41_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,24),
			fetch              => s_fetch(41,24),
			data_in            => s_data_in(41,24),
			data_out           => s_data_out(41,24),
			out1               => s_out1(41,24),
			out2               => s_out2(41,24),
			lock_lower_row_out => s_locks_lower_out(41,24),
			lock_lower_row_in  => s_locks_lower_in(41,24),
			in1                => s_in1(41,24),
			in2                => s_in2(41,24),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(24)
		);
	s_in1(41,24)            <= s_out1(42,24);
	s_in2(41,24)            <= s_out2(42,25);
	s_locks_lower_in(41,24) <= s_locks_lower_out(42,24);

		normal_cell_41_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,25),
			fetch              => s_fetch(41,25),
			data_in            => s_data_in(41,25),
			data_out           => s_data_out(41,25),
			out1               => s_out1(41,25),
			out2               => s_out2(41,25),
			lock_lower_row_out => s_locks_lower_out(41,25),
			lock_lower_row_in  => s_locks_lower_in(41,25),
			in1                => s_in1(41,25),
			in2                => s_in2(41,25),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(25)
		);
	s_in1(41,25)            <= s_out1(42,25);
	s_in2(41,25)            <= s_out2(42,26);
	s_locks_lower_in(41,25) <= s_locks_lower_out(42,25);

		normal_cell_41_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,26),
			fetch              => s_fetch(41,26),
			data_in            => s_data_in(41,26),
			data_out           => s_data_out(41,26),
			out1               => s_out1(41,26),
			out2               => s_out2(41,26),
			lock_lower_row_out => s_locks_lower_out(41,26),
			lock_lower_row_in  => s_locks_lower_in(41,26),
			in1                => s_in1(41,26),
			in2                => s_in2(41,26),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(26)
		);
	s_in1(41,26)            <= s_out1(42,26);
	s_in2(41,26)            <= s_out2(42,27);
	s_locks_lower_in(41,26) <= s_locks_lower_out(42,26);

		normal_cell_41_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,27),
			fetch              => s_fetch(41,27),
			data_in            => s_data_in(41,27),
			data_out           => s_data_out(41,27),
			out1               => s_out1(41,27),
			out2               => s_out2(41,27),
			lock_lower_row_out => s_locks_lower_out(41,27),
			lock_lower_row_in  => s_locks_lower_in(41,27),
			in1                => s_in1(41,27),
			in2                => s_in2(41,27),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(27)
		);
	s_in1(41,27)            <= s_out1(42,27);
	s_in2(41,27)            <= s_out2(42,28);
	s_locks_lower_in(41,27) <= s_locks_lower_out(42,27);

		normal_cell_41_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,28),
			fetch              => s_fetch(41,28),
			data_in            => s_data_in(41,28),
			data_out           => s_data_out(41,28),
			out1               => s_out1(41,28),
			out2               => s_out2(41,28),
			lock_lower_row_out => s_locks_lower_out(41,28),
			lock_lower_row_in  => s_locks_lower_in(41,28),
			in1                => s_in1(41,28),
			in2                => s_in2(41,28),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(28)
		);
	s_in1(41,28)            <= s_out1(42,28);
	s_in2(41,28)            <= s_out2(42,29);
	s_locks_lower_in(41,28) <= s_locks_lower_out(42,28);

		normal_cell_41_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,29),
			fetch              => s_fetch(41,29),
			data_in            => s_data_in(41,29),
			data_out           => s_data_out(41,29),
			out1               => s_out1(41,29),
			out2               => s_out2(41,29),
			lock_lower_row_out => s_locks_lower_out(41,29),
			lock_lower_row_in  => s_locks_lower_in(41,29),
			in1                => s_in1(41,29),
			in2                => s_in2(41,29),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(29)
		);
	s_in1(41,29)            <= s_out1(42,29);
	s_in2(41,29)            <= s_out2(42,30);
	s_locks_lower_in(41,29) <= s_locks_lower_out(42,29);

		normal_cell_41_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,30),
			fetch              => s_fetch(41,30),
			data_in            => s_data_in(41,30),
			data_out           => s_data_out(41,30),
			out1               => s_out1(41,30),
			out2               => s_out2(41,30),
			lock_lower_row_out => s_locks_lower_out(41,30),
			lock_lower_row_in  => s_locks_lower_in(41,30),
			in1                => s_in1(41,30),
			in2                => s_in2(41,30),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(30)
		);
	s_in1(41,30)            <= s_out1(42,30);
	s_in2(41,30)            <= s_out2(42,31);
	s_locks_lower_in(41,30) <= s_locks_lower_out(42,30);

		normal_cell_41_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,31),
			fetch              => s_fetch(41,31),
			data_in            => s_data_in(41,31),
			data_out           => s_data_out(41,31),
			out1               => s_out1(41,31),
			out2               => s_out2(41,31),
			lock_lower_row_out => s_locks_lower_out(41,31),
			lock_lower_row_in  => s_locks_lower_in(41,31),
			in1                => s_in1(41,31),
			in2                => s_in2(41,31),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(31)
		);
	s_in1(41,31)            <= s_out1(42,31);
	s_in2(41,31)            <= s_out2(42,32);
	s_locks_lower_in(41,31) <= s_locks_lower_out(42,31);

		normal_cell_41_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,32),
			fetch              => s_fetch(41,32),
			data_in            => s_data_in(41,32),
			data_out           => s_data_out(41,32),
			out1               => s_out1(41,32),
			out2               => s_out2(41,32),
			lock_lower_row_out => s_locks_lower_out(41,32),
			lock_lower_row_in  => s_locks_lower_in(41,32),
			in1                => s_in1(41,32),
			in2                => s_in2(41,32),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(32)
		);
	s_in1(41,32)            <= s_out1(42,32);
	s_in2(41,32)            <= s_out2(42,33);
	s_locks_lower_in(41,32) <= s_locks_lower_out(42,32);

		normal_cell_41_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,33),
			fetch              => s_fetch(41,33),
			data_in            => s_data_in(41,33),
			data_out           => s_data_out(41,33),
			out1               => s_out1(41,33),
			out2               => s_out2(41,33),
			lock_lower_row_out => s_locks_lower_out(41,33),
			lock_lower_row_in  => s_locks_lower_in(41,33),
			in1                => s_in1(41,33),
			in2                => s_in2(41,33),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(33)
		);
	s_in1(41,33)            <= s_out1(42,33);
	s_in2(41,33)            <= s_out2(42,34);
	s_locks_lower_in(41,33) <= s_locks_lower_out(42,33);

		normal_cell_41_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,34),
			fetch              => s_fetch(41,34),
			data_in            => s_data_in(41,34),
			data_out           => s_data_out(41,34),
			out1               => s_out1(41,34),
			out2               => s_out2(41,34),
			lock_lower_row_out => s_locks_lower_out(41,34),
			lock_lower_row_in  => s_locks_lower_in(41,34),
			in1                => s_in1(41,34),
			in2                => s_in2(41,34),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(34)
		);
	s_in1(41,34)            <= s_out1(42,34);
	s_in2(41,34)            <= s_out2(42,35);
	s_locks_lower_in(41,34) <= s_locks_lower_out(42,34);

		normal_cell_41_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,35),
			fetch              => s_fetch(41,35),
			data_in            => s_data_in(41,35),
			data_out           => s_data_out(41,35),
			out1               => s_out1(41,35),
			out2               => s_out2(41,35),
			lock_lower_row_out => s_locks_lower_out(41,35),
			lock_lower_row_in  => s_locks_lower_in(41,35),
			in1                => s_in1(41,35),
			in2                => s_in2(41,35),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(35)
		);
	s_in1(41,35)            <= s_out1(42,35);
	s_in2(41,35)            <= s_out2(42,36);
	s_locks_lower_in(41,35) <= s_locks_lower_out(42,35);

		normal_cell_41_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,36),
			fetch              => s_fetch(41,36),
			data_in            => s_data_in(41,36),
			data_out           => s_data_out(41,36),
			out1               => s_out1(41,36),
			out2               => s_out2(41,36),
			lock_lower_row_out => s_locks_lower_out(41,36),
			lock_lower_row_in  => s_locks_lower_in(41,36),
			in1                => s_in1(41,36),
			in2                => s_in2(41,36),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(36)
		);
	s_in1(41,36)            <= s_out1(42,36);
	s_in2(41,36)            <= s_out2(42,37);
	s_locks_lower_in(41,36) <= s_locks_lower_out(42,36);

		normal_cell_41_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,37),
			fetch              => s_fetch(41,37),
			data_in            => s_data_in(41,37),
			data_out           => s_data_out(41,37),
			out1               => s_out1(41,37),
			out2               => s_out2(41,37),
			lock_lower_row_out => s_locks_lower_out(41,37),
			lock_lower_row_in  => s_locks_lower_in(41,37),
			in1                => s_in1(41,37),
			in2                => s_in2(41,37),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(37)
		);
	s_in1(41,37)            <= s_out1(42,37);
	s_in2(41,37)            <= s_out2(42,38);
	s_locks_lower_in(41,37) <= s_locks_lower_out(42,37);

		normal_cell_41_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,38),
			fetch              => s_fetch(41,38),
			data_in            => s_data_in(41,38),
			data_out           => s_data_out(41,38),
			out1               => s_out1(41,38),
			out2               => s_out2(41,38),
			lock_lower_row_out => s_locks_lower_out(41,38),
			lock_lower_row_in  => s_locks_lower_in(41,38),
			in1                => s_in1(41,38),
			in2                => s_in2(41,38),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(38)
		);
	s_in1(41,38)            <= s_out1(42,38);
	s_in2(41,38)            <= s_out2(42,39);
	s_locks_lower_in(41,38) <= s_locks_lower_out(42,38);

		normal_cell_41_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,39),
			fetch              => s_fetch(41,39),
			data_in            => s_data_in(41,39),
			data_out           => s_data_out(41,39),
			out1               => s_out1(41,39),
			out2               => s_out2(41,39),
			lock_lower_row_out => s_locks_lower_out(41,39),
			lock_lower_row_in  => s_locks_lower_in(41,39),
			in1                => s_in1(41,39),
			in2                => s_in2(41,39),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(39)
		);
	s_in1(41,39)            <= s_out1(42,39);
	s_in2(41,39)            <= s_out2(42,40);
	s_locks_lower_in(41,39) <= s_locks_lower_out(42,39);

		normal_cell_41_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,40),
			fetch              => s_fetch(41,40),
			data_in            => s_data_in(41,40),
			data_out           => s_data_out(41,40),
			out1               => s_out1(41,40),
			out2               => s_out2(41,40),
			lock_lower_row_out => s_locks_lower_out(41,40),
			lock_lower_row_in  => s_locks_lower_in(41,40),
			in1                => s_in1(41,40),
			in2                => s_in2(41,40),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(40)
		);
	s_in1(41,40)            <= s_out1(42,40);
	s_in2(41,40)            <= s_out2(42,41);
	s_locks_lower_in(41,40) <= s_locks_lower_out(42,40);

		normal_cell_41_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,41),
			fetch              => s_fetch(41,41),
			data_in            => s_data_in(41,41),
			data_out           => s_data_out(41,41),
			out1               => s_out1(41,41),
			out2               => s_out2(41,41),
			lock_lower_row_out => s_locks_lower_out(41,41),
			lock_lower_row_in  => s_locks_lower_in(41,41),
			in1                => s_in1(41,41),
			in2                => s_in2(41,41),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(41)
		);
	s_in1(41,41)            <= s_out1(42,41);
	s_in2(41,41)            <= s_out2(42,42);
	s_locks_lower_in(41,41) <= s_locks_lower_out(42,41);

		normal_cell_41_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,42),
			fetch              => s_fetch(41,42),
			data_in            => s_data_in(41,42),
			data_out           => s_data_out(41,42),
			out1               => s_out1(41,42),
			out2               => s_out2(41,42),
			lock_lower_row_out => s_locks_lower_out(41,42),
			lock_lower_row_in  => s_locks_lower_in(41,42),
			in1                => s_in1(41,42),
			in2                => s_in2(41,42),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(42)
		);
	s_in1(41,42)            <= s_out1(42,42);
	s_in2(41,42)            <= s_out2(42,43);
	s_locks_lower_in(41,42) <= s_locks_lower_out(42,42);

		normal_cell_41_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,43),
			fetch              => s_fetch(41,43),
			data_in            => s_data_in(41,43),
			data_out           => s_data_out(41,43),
			out1               => s_out1(41,43),
			out2               => s_out2(41,43),
			lock_lower_row_out => s_locks_lower_out(41,43),
			lock_lower_row_in  => s_locks_lower_in(41,43),
			in1                => s_in1(41,43),
			in2                => s_in2(41,43),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(43)
		);
	s_in1(41,43)            <= s_out1(42,43);
	s_in2(41,43)            <= s_out2(42,44);
	s_locks_lower_in(41,43) <= s_locks_lower_out(42,43);

		normal_cell_41_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,44),
			fetch              => s_fetch(41,44),
			data_in            => s_data_in(41,44),
			data_out           => s_data_out(41,44),
			out1               => s_out1(41,44),
			out2               => s_out2(41,44),
			lock_lower_row_out => s_locks_lower_out(41,44),
			lock_lower_row_in  => s_locks_lower_in(41,44),
			in1                => s_in1(41,44),
			in2                => s_in2(41,44),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(44)
		);
	s_in1(41,44)            <= s_out1(42,44);
	s_in2(41,44)            <= s_out2(42,45);
	s_locks_lower_in(41,44) <= s_locks_lower_out(42,44);

		normal_cell_41_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,45),
			fetch              => s_fetch(41,45),
			data_in            => s_data_in(41,45),
			data_out           => s_data_out(41,45),
			out1               => s_out1(41,45),
			out2               => s_out2(41,45),
			lock_lower_row_out => s_locks_lower_out(41,45),
			lock_lower_row_in  => s_locks_lower_in(41,45),
			in1                => s_in1(41,45),
			in2                => s_in2(41,45),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(45)
		);
	s_in1(41,45)            <= s_out1(42,45);
	s_in2(41,45)            <= s_out2(42,46);
	s_locks_lower_in(41,45) <= s_locks_lower_out(42,45);

		normal_cell_41_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,46),
			fetch              => s_fetch(41,46),
			data_in            => s_data_in(41,46),
			data_out           => s_data_out(41,46),
			out1               => s_out1(41,46),
			out2               => s_out2(41,46),
			lock_lower_row_out => s_locks_lower_out(41,46),
			lock_lower_row_in  => s_locks_lower_in(41,46),
			in1                => s_in1(41,46),
			in2                => s_in2(41,46),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(46)
		);
	s_in1(41,46)            <= s_out1(42,46);
	s_in2(41,46)            <= s_out2(42,47);
	s_locks_lower_in(41,46) <= s_locks_lower_out(42,46);

		normal_cell_41_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,47),
			fetch              => s_fetch(41,47),
			data_in            => s_data_in(41,47),
			data_out           => s_data_out(41,47),
			out1               => s_out1(41,47),
			out2               => s_out2(41,47),
			lock_lower_row_out => s_locks_lower_out(41,47),
			lock_lower_row_in  => s_locks_lower_in(41,47),
			in1                => s_in1(41,47),
			in2                => s_in2(41,47),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(47)
		);
	s_in1(41,47)            <= s_out1(42,47);
	s_in2(41,47)            <= s_out2(42,48);
	s_locks_lower_in(41,47) <= s_locks_lower_out(42,47);

		normal_cell_41_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,48),
			fetch              => s_fetch(41,48),
			data_in            => s_data_in(41,48),
			data_out           => s_data_out(41,48),
			out1               => s_out1(41,48),
			out2               => s_out2(41,48),
			lock_lower_row_out => s_locks_lower_out(41,48),
			lock_lower_row_in  => s_locks_lower_in(41,48),
			in1                => s_in1(41,48),
			in2                => s_in2(41,48),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(48)
		);
	s_in1(41,48)            <= s_out1(42,48);
	s_in2(41,48)            <= s_out2(42,49);
	s_locks_lower_in(41,48) <= s_locks_lower_out(42,48);

		normal_cell_41_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,49),
			fetch              => s_fetch(41,49),
			data_in            => s_data_in(41,49),
			data_out           => s_data_out(41,49),
			out1               => s_out1(41,49),
			out2               => s_out2(41,49),
			lock_lower_row_out => s_locks_lower_out(41,49),
			lock_lower_row_in  => s_locks_lower_in(41,49),
			in1                => s_in1(41,49),
			in2                => s_in2(41,49),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(49)
		);
	s_in1(41,49)            <= s_out1(42,49);
	s_in2(41,49)            <= s_out2(42,50);
	s_locks_lower_in(41,49) <= s_locks_lower_out(42,49);

		normal_cell_41_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,50),
			fetch              => s_fetch(41,50),
			data_in            => s_data_in(41,50),
			data_out           => s_data_out(41,50),
			out1               => s_out1(41,50),
			out2               => s_out2(41,50),
			lock_lower_row_out => s_locks_lower_out(41,50),
			lock_lower_row_in  => s_locks_lower_in(41,50),
			in1                => s_in1(41,50),
			in2                => s_in2(41,50),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(50)
		);
	s_in1(41,50)            <= s_out1(42,50);
	s_in2(41,50)            <= s_out2(42,51);
	s_locks_lower_in(41,50) <= s_locks_lower_out(42,50);

		normal_cell_41_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,51),
			fetch              => s_fetch(41,51),
			data_in            => s_data_in(41,51),
			data_out           => s_data_out(41,51),
			out1               => s_out1(41,51),
			out2               => s_out2(41,51),
			lock_lower_row_out => s_locks_lower_out(41,51),
			lock_lower_row_in  => s_locks_lower_in(41,51),
			in1                => s_in1(41,51),
			in2                => s_in2(41,51),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(51)
		);
	s_in1(41,51)            <= s_out1(42,51);
	s_in2(41,51)            <= s_out2(42,52);
	s_locks_lower_in(41,51) <= s_locks_lower_out(42,51);

		normal_cell_41_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,52),
			fetch              => s_fetch(41,52),
			data_in            => s_data_in(41,52),
			data_out           => s_data_out(41,52),
			out1               => s_out1(41,52),
			out2               => s_out2(41,52),
			lock_lower_row_out => s_locks_lower_out(41,52),
			lock_lower_row_in  => s_locks_lower_in(41,52),
			in1                => s_in1(41,52),
			in2                => s_in2(41,52),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(52)
		);
	s_in1(41,52)            <= s_out1(42,52);
	s_in2(41,52)            <= s_out2(42,53);
	s_locks_lower_in(41,52) <= s_locks_lower_out(42,52);

		normal_cell_41_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,53),
			fetch              => s_fetch(41,53),
			data_in            => s_data_in(41,53),
			data_out           => s_data_out(41,53),
			out1               => s_out1(41,53),
			out2               => s_out2(41,53),
			lock_lower_row_out => s_locks_lower_out(41,53),
			lock_lower_row_in  => s_locks_lower_in(41,53),
			in1                => s_in1(41,53),
			in2                => s_in2(41,53),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(53)
		);
	s_in1(41,53)            <= s_out1(42,53);
	s_in2(41,53)            <= s_out2(42,54);
	s_locks_lower_in(41,53) <= s_locks_lower_out(42,53);

		normal_cell_41_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,54),
			fetch              => s_fetch(41,54),
			data_in            => s_data_in(41,54),
			data_out           => s_data_out(41,54),
			out1               => s_out1(41,54),
			out2               => s_out2(41,54),
			lock_lower_row_out => s_locks_lower_out(41,54),
			lock_lower_row_in  => s_locks_lower_in(41,54),
			in1                => s_in1(41,54),
			in2                => s_in2(41,54),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(54)
		);
	s_in1(41,54)            <= s_out1(42,54);
	s_in2(41,54)            <= s_out2(42,55);
	s_locks_lower_in(41,54) <= s_locks_lower_out(42,54);

		normal_cell_41_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,55),
			fetch              => s_fetch(41,55),
			data_in            => s_data_in(41,55),
			data_out           => s_data_out(41,55),
			out1               => s_out1(41,55),
			out2               => s_out2(41,55),
			lock_lower_row_out => s_locks_lower_out(41,55),
			lock_lower_row_in  => s_locks_lower_in(41,55),
			in1                => s_in1(41,55),
			in2                => s_in2(41,55),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(55)
		);
	s_in1(41,55)            <= s_out1(42,55);
	s_in2(41,55)            <= s_out2(42,56);
	s_locks_lower_in(41,55) <= s_locks_lower_out(42,55);

		normal_cell_41_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,56),
			fetch              => s_fetch(41,56),
			data_in            => s_data_in(41,56),
			data_out           => s_data_out(41,56),
			out1               => s_out1(41,56),
			out2               => s_out2(41,56),
			lock_lower_row_out => s_locks_lower_out(41,56),
			lock_lower_row_in  => s_locks_lower_in(41,56),
			in1                => s_in1(41,56),
			in2                => s_in2(41,56),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(56)
		);
	s_in1(41,56)            <= s_out1(42,56);
	s_in2(41,56)            <= s_out2(42,57);
	s_locks_lower_in(41,56) <= s_locks_lower_out(42,56);

		normal_cell_41_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,57),
			fetch              => s_fetch(41,57),
			data_in            => s_data_in(41,57),
			data_out           => s_data_out(41,57),
			out1               => s_out1(41,57),
			out2               => s_out2(41,57),
			lock_lower_row_out => s_locks_lower_out(41,57),
			lock_lower_row_in  => s_locks_lower_in(41,57),
			in1                => s_in1(41,57),
			in2                => s_in2(41,57),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(57)
		);
	s_in1(41,57)            <= s_out1(42,57);
	s_in2(41,57)            <= s_out2(42,58);
	s_locks_lower_in(41,57) <= s_locks_lower_out(42,57);

		normal_cell_41_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,58),
			fetch              => s_fetch(41,58),
			data_in            => s_data_in(41,58),
			data_out           => s_data_out(41,58),
			out1               => s_out1(41,58),
			out2               => s_out2(41,58),
			lock_lower_row_out => s_locks_lower_out(41,58),
			lock_lower_row_in  => s_locks_lower_in(41,58),
			in1                => s_in1(41,58),
			in2                => s_in2(41,58),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(58)
		);
	s_in1(41,58)            <= s_out1(42,58);
	s_in2(41,58)            <= s_out2(42,59);
	s_locks_lower_in(41,58) <= s_locks_lower_out(42,58);

		normal_cell_41_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,59),
			fetch              => s_fetch(41,59),
			data_in            => s_data_in(41,59),
			data_out           => s_data_out(41,59),
			out1               => s_out1(41,59),
			out2               => s_out2(41,59),
			lock_lower_row_out => s_locks_lower_out(41,59),
			lock_lower_row_in  => s_locks_lower_in(41,59),
			in1                => s_in1(41,59),
			in2                => s_in2(41,59),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(59)
		);
	s_in1(41,59)            <= s_out1(42,59);
	s_in2(41,59)            <= s_out2(42,60);
	s_locks_lower_in(41,59) <= s_locks_lower_out(42,59);

		last_col_cell_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(41,60),
			fetch              => s_fetch(41,60),
			data_in            => s_data_in(41,60),
			data_out           => s_data_out(41,60),
			out1               => s_out1(41,60),
			out2               => s_out2(41,60),
			lock_lower_row_out => s_locks_lower_out(41,60),
			lock_lower_row_in  => s_locks_lower_in(41,60),
			in1                => s_in1(41,60),
			in2                => (others => '0'),
			lock_row           => s_locks(41),
			piv_found          => s_piv_found,
			row_data           => s_row_data(41),
			col_data           => s_col_data(60)
		);
	s_in1(41,60)            <= s_out1(42,60);
	s_locks_lower_in(41,60) <= s_locks_lower_out(42,60);

		normal_cell_42_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,1),
			fetch              => s_fetch(42,1),
			data_in            => s_data_in(42,1),
			data_out           => s_data_out(42,1),
			out1               => s_out1(42,1),
			out2               => s_out2(42,1),
			lock_lower_row_out => s_locks_lower_out(42,1),
			lock_lower_row_in  => s_locks_lower_in(42,1),
			in1                => s_in1(42,1),
			in2                => s_in2(42,1),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(1)
		);
	s_in1(42,1)            <= s_out1(43,1);
	s_in2(42,1)            <= s_out2(43,2);
	s_locks_lower_in(42,1) <= s_locks_lower_out(43,1);

		normal_cell_42_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,2),
			fetch              => s_fetch(42,2),
			data_in            => s_data_in(42,2),
			data_out           => s_data_out(42,2),
			out1               => s_out1(42,2),
			out2               => s_out2(42,2),
			lock_lower_row_out => s_locks_lower_out(42,2),
			lock_lower_row_in  => s_locks_lower_in(42,2),
			in1                => s_in1(42,2),
			in2                => s_in2(42,2),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(2)
		);
	s_in1(42,2)            <= s_out1(43,2);
	s_in2(42,2)            <= s_out2(43,3);
	s_locks_lower_in(42,2) <= s_locks_lower_out(43,2);

		normal_cell_42_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,3),
			fetch              => s_fetch(42,3),
			data_in            => s_data_in(42,3),
			data_out           => s_data_out(42,3),
			out1               => s_out1(42,3),
			out2               => s_out2(42,3),
			lock_lower_row_out => s_locks_lower_out(42,3),
			lock_lower_row_in  => s_locks_lower_in(42,3),
			in1                => s_in1(42,3),
			in2                => s_in2(42,3),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(3)
		);
	s_in1(42,3)            <= s_out1(43,3);
	s_in2(42,3)            <= s_out2(43,4);
	s_locks_lower_in(42,3) <= s_locks_lower_out(43,3);

		normal_cell_42_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,4),
			fetch              => s_fetch(42,4),
			data_in            => s_data_in(42,4),
			data_out           => s_data_out(42,4),
			out1               => s_out1(42,4),
			out2               => s_out2(42,4),
			lock_lower_row_out => s_locks_lower_out(42,4),
			lock_lower_row_in  => s_locks_lower_in(42,4),
			in1                => s_in1(42,4),
			in2                => s_in2(42,4),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(4)
		);
	s_in1(42,4)            <= s_out1(43,4);
	s_in2(42,4)            <= s_out2(43,5);
	s_locks_lower_in(42,4) <= s_locks_lower_out(43,4);

		normal_cell_42_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,5),
			fetch              => s_fetch(42,5),
			data_in            => s_data_in(42,5),
			data_out           => s_data_out(42,5),
			out1               => s_out1(42,5),
			out2               => s_out2(42,5),
			lock_lower_row_out => s_locks_lower_out(42,5),
			lock_lower_row_in  => s_locks_lower_in(42,5),
			in1                => s_in1(42,5),
			in2                => s_in2(42,5),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(5)
		);
	s_in1(42,5)            <= s_out1(43,5);
	s_in2(42,5)            <= s_out2(43,6);
	s_locks_lower_in(42,5) <= s_locks_lower_out(43,5);

		normal_cell_42_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,6),
			fetch              => s_fetch(42,6),
			data_in            => s_data_in(42,6),
			data_out           => s_data_out(42,6),
			out1               => s_out1(42,6),
			out2               => s_out2(42,6),
			lock_lower_row_out => s_locks_lower_out(42,6),
			lock_lower_row_in  => s_locks_lower_in(42,6),
			in1                => s_in1(42,6),
			in2                => s_in2(42,6),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(6)
		);
	s_in1(42,6)            <= s_out1(43,6);
	s_in2(42,6)            <= s_out2(43,7);
	s_locks_lower_in(42,6) <= s_locks_lower_out(43,6);

		normal_cell_42_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,7),
			fetch              => s_fetch(42,7),
			data_in            => s_data_in(42,7),
			data_out           => s_data_out(42,7),
			out1               => s_out1(42,7),
			out2               => s_out2(42,7),
			lock_lower_row_out => s_locks_lower_out(42,7),
			lock_lower_row_in  => s_locks_lower_in(42,7),
			in1                => s_in1(42,7),
			in2                => s_in2(42,7),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(7)
		);
	s_in1(42,7)            <= s_out1(43,7);
	s_in2(42,7)            <= s_out2(43,8);
	s_locks_lower_in(42,7) <= s_locks_lower_out(43,7);

		normal_cell_42_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,8),
			fetch              => s_fetch(42,8),
			data_in            => s_data_in(42,8),
			data_out           => s_data_out(42,8),
			out1               => s_out1(42,8),
			out2               => s_out2(42,8),
			lock_lower_row_out => s_locks_lower_out(42,8),
			lock_lower_row_in  => s_locks_lower_in(42,8),
			in1                => s_in1(42,8),
			in2                => s_in2(42,8),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(8)
		);
	s_in1(42,8)            <= s_out1(43,8);
	s_in2(42,8)            <= s_out2(43,9);
	s_locks_lower_in(42,8) <= s_locks_lower_out(43,8);

		normal_cell_42_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,9),
			fetch              => s_fetch(42,9),
			data_in            => s_data_in(42,9),
			data_out           => s_data_out(42,9),
			out1               => s_out1(42,9),
			out2               => s_out2(42,9),
			lock_lower_row_out => s_locks_lower_out(42,9),
			lock_lower_row_in  => s_locks_lower_in(42,9),
			in1                => s_in1(42,9),
			in2                => s_in2(42,9),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(9)
		);
	s_in1(42,9)            <= s_out1(43,9);
	s_in2(42,9)            <= s_out2(43,10);
	s_locks_lower_in(42,9) <= s_locks_lower_out(43,9);

		normal_cell_42_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,10),
			fetch              => s_fetch(42,10),
			data_in            => s_data_in(42,10),
			data_out           => s_data_out(42,10),
			out1               => s_out1(42,10),
			out2               => s_out2(42,10),
			lock_lower_row_out => s_locks_lower_out(42,10),
			lock_lower_row_in  => s_locks_lower_in(42,10),
			in1                => s_in1(42,10),
			in2                => s_in2(42,10),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(10)
		);
	s_in1(42,10)            <= s_out1(43,10);
	s_in2(42,10)            <= s_out2(43,11);
	s_locks_lower_in(42,10) <= s_locks_lower_out(43,10);

		normal_cell_42_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,11),
			fetch              => s_fetch(42,11),
			data_in            => s_data_in(42,11),
			data_out           => s_data_out(42,11),
			out1               => s_out1(42,11),
			out2               => s_out2(42,11),
			lock_lower_row_out => s_locks_lower_out(42,11),
			lock_lower_row_in  => s_locks_lower_in(42,11),
			in1                => s_in1(42,11),
			in2                => s_in2(42,11),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(11)
		);
	s_in1(42,11)            <= s_out1(43,11);
	s_in2(42,11)            <= s_out2(43,12);
	s_locks_lower_in(42,11) <= s_locks_lower_out(43,11);

		normal_cell_42_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,12),
			fetch              => s_fetch(42,12),
			data_in            => s_data_in(42,12),
			data_out           => s_data_out(42,12),
			out1               => s_out1(42,12),
			out2               => s_out2(42,12),
			lock_lower_row_out => s_locks_lower_out(42,12),
			lock_lower_row_in  => s_locks_lower_in(42,12),
			in1                => s_in1(42,12),
			in2                => s_in2(42,12),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(12)
		);
	s_in1(42,12)            <= s_out1(43,12);
	s_in2(42,12)            <= s_out2(43,13);
	s_locks_lower_in(42,12) <= s_locks_lower_out(43,12);

		normal_cell_42_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,13),
			fetch              => s_fetch(42,13),
			data_in            => s_data_in(42,13),
			data_out           => s_data_out(42,13),
			out1               => s_out1(42,13),
			out2               => s_out2(42,13),
			lock_lower_row_out => s_locks_lower_out(42,13),
			lock_lower_row_in  => s_locks_lower_in(42,13),
			in1                => s_in1(42,13),
			in2                => s_in2(42,13),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(13)
		);
	s_in1(42,13)            <= s_out1(43,13);
	s_in2(42,13)            <= s_out2(43,14);
	s_locks_lower_in(42,13) <= s_locks_lower_out(43,13);

		normal_cell_42_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,14),
			fetch              => s_fetch(42,14),
			data_in            => s_data_in(42,14),
			data_out           => s_data_out(42,14),
			out1               => s_out1(42,14),
			out2               => s_out2(42,14),
			lock_lower_row_out => s_locks_lower_out(42,14),
			lock_lower_row_in  => s_locks_lower_in(42,14),
			in1                => s_in1(42,14),
			in2                => s_in2(42,14),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(14)
		);
	s_in1(42,14)            <= s_out1(43,14);
	s_in2(42,14)            <= s_out2(43,15);
	s_locks_lower_in(42,14) <= s_locks_lower_out(43,14);

		normal_cell_42_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,15),
			fetch              => s_fetch(42,15),
			data_in            => s_data_in(42,15),
			data_out           => s_data_out(42,15),
			out1               => s_out1(42,15),
			out2               => s_out2(42,15),
			lock_lower_row_out => s_locks_lower_out(42,15),
			lock_lower_row_in  => s_locks_lower_in(42,15),
			in1                => s_in1(42,15),
			in2                => s_in2(42,15),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(15)
		);
	s_in1(42,15)            <= s_out1(43,15);
	s_in2(42,15)            <= s_out2(43,16);
	s_locks_lower_in(42,15) <= s_locks_lower_out(43,15);

		normal_cell_42_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,16),
			fetch              => s_fetch(42,16),
			data_in            => s_data_in(42,16),
			data_out           => s_data_out(42,16),
			out1               => s_out1(42,16),
			out2               => s_out2(42,16),
			lock_lower_row_out => s_locks_lower_out(42,16),
			lock_lower_row_in  => s_locks_lower_in(42,16),
			in1                => s_in1(42,16),
			in2                => s_in2(42,16),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(16)
		);
	s_in1(42,16)            <= s_out1(43,16);
	s_in2(42,16)            <= s_out2(43,17);
	s_locks_lower_in(42,16) <= s_locks_lower_out(43,16);

		normal_cell_42_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,17),
			fetch              => s_fetch(42,17),
			data_in            => s_data_in(42,17),
			data_out           => s_data_out(42,17),
			out1               => s_out1(42,17),
			out2               => s_out2(42,17),
			lock_lower_row_out => s_locks_lower_out(42,17),
			lock_lower_row_in  => s_locks_lower_in(42,17),
			in1                => s_in1(42,17),
			in2                => s_in2(42,17),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(17)
		);
	s_in1(42,17)            <= s_out1(43,17);
	s_in2(42,17)            <= s_out2(43,18);
	s_locks_lower_in(42,17) <= s_locks_lower_out(43,17);

		normal_cell_42_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,18),
			fetch              => s_fetch(42,18),
			data_in            => s_data_in(42,18),
			data_out           => s_data_out(42,18),
			out1               => s_out1(42,18),
			out2               => s_out2(42,18),
			lock_lower_row_out => s_locks_lower_out(42,18),
			lock_lower_row_in  => s_locks_lower_in(42,18),
			in1                => s_in1(42,18),
			in2                => s_in2(42,18),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(18)
		);
	s_in1(42,18)            <= s_out1(43,18);
	s_in2(42,18)            <= s_out2(43,19);
	s_locks_lower_in(42,18) <= s_locks_lower_out(43,18);

		normal_cell_42_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,19),
			fetch              => s_fetch(42,19),
			data_in            => s_data_in(42,19),
			data_out           => s_data_out(42,19),
			out1               => s_out1(42,19),
			out2               => s_out2(42,19),
			lock_lower_row_out => s_locks_lower_out(42,19),
			lock_lower_row_in  => s_locks_lower_in(42,19),
			in1                => s_in1(42,19),
			in2                => s_in2(42,19),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(19)
		);
	s_in1(42,19)            <= s_out1(43,19);
	s_in2(42,19)            <= s_out2(43,20);
	s_locks_lower_in(42,19) <= s_locks_lower_out(43,19);

		normal_cell_42_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,20),
			fetch              => s_fetch(42,20),
			data_in            => s_data_in(42,20),
			data_out           => s_data_out(42,20),
			out1               => s_out1(42,20),
			out2               => s_out2(42,20),
			lock_lower_row_out => s_locks_lower_out(42,20),
			lock_lower_row_in  => s_locks_lower_in(42,20),
			in1                => s_in1(42,20),
			in2                => s_in2(42,20),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(20)
		);
	s_in1(42,20)            <= s_out1(43,20);
	s_in2(42,20)            <= s_out2(43,21);
	s_locks_lower_in(42,20) <= s_locks_lower_out(43,20);

		normal_cell_42_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,21),
			fetch              => s_fetch(42,21),
			data_in            => s_data_in(42,21),
			data_out           => s_data_out(42,21),
			out1               => s_out1(42,21),
			out2               => s_out2(42,21),
			lock_lower_row_out => s_locks_lower_out(42,21),
			lock_lower_row_in  => s_locks_lower_in(42,21),
			in1                => s_in1(42,21),
			in2                => s_in2(42,21),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(21)
		);
	s_in1(42,21)            <= s_out1(43,21);
	s_in2(42,21)            <= s_out2(43,22);
	s_locks_lower_in(42,21) <= s_locks_lower_out(43,21);

		normal_cell_42_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,22),
			fetch              => s_fetch(42,22),
			data_in            => s_data_in(42,22),
			data_out           => s_data_out(42,22),
			out1               => s_out1(42,22),
			out2               => s_out2(42,22),
			lock_lower_row_out => s_locks_lower_out(42,22),
			lock_lower_row_in  => s_locks_lower_in(42,22),
			in1                => s_in1(42,22),
			in2                => s_in2(42,22),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(22)
		);
	s_in1(42,22)            <= s_out1(43,22);
	s_in2(42,22)            <= s_out2(43,23);
	s_locks_lower_in(42,22) <= s_locks_lower_out(43,22);

		normal_cell_42_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,23),
			fetch              => s_fetch(42,23),
			data_in            => s_data_in(42,23),
			data_out           => s_data_out(42,23),
			out1               => s_out1(42,23),
			out2               => s_out2(42,23),
			lock_lower_row_out => s_locks_lower_out(42,23),
			lock_lower_row_in  => s_locks_lower_in(42,23),
			in1                => s_in1(42,23),
			in2                => s_in2(42,23),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(23)
		);
	s_in1(42,23)            <= s_out1(43,23);
	s_in2(42,23)            <= s_out2(43,24);
	s_locks_lower_in(42,23) <= s_locks_lower_out(43,23);

		normal_cell_42_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,24),
			fetch              => s_fetch(42,24),
			data_in            => s_data_in(42,24),
			data_out           => s_data_out(42,24),
			out1               => s_out1(42,24),
			out2               => s_out2(42,24),
			lock_lower_row_out => s_locks_lower_out(42,24),
			lock_lower_row_in  => s_locks_lower_in(42,24),
			in1                => s_in1(42,24),
			in2                => s_in2(42,24),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(24)
		);
	s_in1(42,24)            <= s_out1(43,24);
	s_in2(42,24)            <= s_out2(43,25);
	s_locks_lower_in(42,24) <= s_locks_lower_out(43,24);

		normal_cell_42_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,25),
			fetch              => s_fetch(42,25),
			data_in            => s_data_in(42,25),
			data_out           => s_data_out(42,25),
			out1               => s_out1(42,25),
			out2               => s_out2(42,25),
			lock_lower_row_out => s_locks_lower_out(42,25),
			lock_lower_row_in  => s_locks_lower_in(42,25),
			in1                => s_in1(42,25),
			in2                => s_in2(42,25),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(25)
		);
	s_in1(42,25)            <= s_out1(43,25);
	s_in2(42,25)            <= s_out2(43,26);
	s_locks_lower_in(42,25) <= s_locks_lower_out(43,25);

		normal_cell_42_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,26),
			fetch              => s_fetch(42,26),
			data_in            => s_data_in(42,26),
			data_out           => s_data_out(42,26),
			out1               => s_out1(42,26),
			out2               => s_out2(42,26),
			lock_lower_row_out => s_locks_lower_out(42,26),
			lock_lower_row_in  => s_locks_lower_in(42,26),
			in1                => s_in1(42,26),
			in2                => s_in2(42,26),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(26)
		);
	s_in1(42,26)            <= s_out1(43,26);
	s_in2(42,26)            <= s_out2(43,27);
	s_locks_lower_in(42,26) <= s_locks_lower_out(43,26);

		normal_cell_42_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,27),
			fetch              => s_fetch(42,27),
			data_in            => s_data_in(42,27),
			data_out           => s_data_out(42,27),
			out1               => s_out1(42,27),
			out2               => s_out2(42,27),
			lock_lower_row_out => s_locks_lower_out(42,27),
			lock_lower_row_in  => s_locks_lower_in(42,27),
			in1                => s_in1(42,27),
			in2                => s_in2(42,27),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(27)
		);
	s_in1(42,27)            <= s_out1(43,27);
	s_in2(42,27)            <= s_out2(43,28);
	s_locks_lower_in(42,27) <= s_locks_lower_out(43,27);

		normal_cell_42_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,28),
			fetch              => s_fetch(42,28),
			data_in            => s_data_in(42,28),
			data_out           => s_data_out(42,28),
			out1               => s_out1(42,28),
			out2               => s_out2(42,28),
			lock_lower_row_out => s_locks_lower_out(42,28),
			lock_lower_row_in  => s_locks_lower_in(42,28),
			in1                => s_in1(42,28),
			in2                => s_in2(42,28),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(28)
		);
	s_in1(42,28)            <= s_out1(43,28);
	s_in2(42,28)            <= s_out2(43,29);
	s_locks_lower_in(42,28) <= s_locks_lower_out(43,28);

		normal_cell_42_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,29),
			fetch              => s_fetch(42,29),
			data_in            => s_data_in(42,29),
			data_out           => s_data_out(42,29),
			out1               => s_out1(42,29),
			out2               => s_out2(42,29),
			lock_lower_row_out => s_locks_lower_out(42,29),
			lock_lower_row_in  => s_locks_lower_in(42,29),
			in1                => s_in1(42,29),
			in2                => s_in2(42,29),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(29)
		);
	s_in1(42,29)            <= s_out1(43,29);
	s_in2(42,29)            <= s_out2(43,30);
	s_locks_lower_in(42,29) <= s_locks_lower_out(43,29);

		normal_cell_42_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,30),
			fetch              => s_fetch(42,30),
			data_in            => s_data_in(42,30),
			data_out           => s_data_out(42,30),
			out1               => s_out1(42,30),
			out2               => s_out2(42,30),
			lock_lower_row_out => s_locks_lower_out(42,30),
			lock_lower_row_in  => s_locks_lower_in(42,30),
			in1                => s_in1(42,30),
			in2                => s_in2(42,30),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(30)
		);
	s_in1(42,30)            <= s_out1(43,30);
	s_in2(42,30)            <= s_out2(43,31);
	s_locks_lower_in(42,30) <= s_locks_lower_out(43,30);

		normal_cell_42_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,31),
			fetch              => s_fetch(42,31),
			data_in            => s_data_in(42,31),
			data_out           => s_data_out(42,31),
			out1               => s_out1(42,31),
			out2               => s_out2(42,31),
			lock_lower_row_out => s_locks_lower_out(42,31),
			lock_lower_row_in  => s_locks_lower_in(42,31),
			in1                => s_in1(42,31),
			in2                => s_in2(42,31),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(31)
		);
	s_in1(42,31)            <= s_out1(43,31);
	s_in2(42,31)            <= s_out2(43,32);
	s_locks_lower_in(42,31) <= s_locks_lower_out(43,31);

		normal_cell_42_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,32),
			fetch              => s_fetch(42,32),
			data_in            => s_data_in(42,32),
			data_out           => s_data_out(42,32),
			out1               => s_out1(42,32),
			out2               => s_out2(42,32),
			lock_lower_row_out => s_locks_lower_out(42,32),
			lock_lower_row_in  => s_locks_lower_in(42,32),
			in1                => s_in1(42,32),
			in2                => s_in2(42,32),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(32)
		);
	s_in1(42,32)            <= s_out1(43,32);
	s_in2(42,32)            <= s_out2(43,33);
	s_locks_lower_in(42,32) <= s_locks_lower_out(43,32);

		normal_cell_42_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,33),
			fetch              => s_fetch(42,33),
			data_in            => s_data_in(42,33),
			data_out           => s_data_out(42,33),
			out1               => s_out1(42,33),
			out2               => s_out2(42,33),
			lock_lower_row_out => s_locks_lower_out(42,33),
			lock_lower_row_in  => s_locks_lower_in(42,33),
			in1                => s_in1(42,33),
			in2                => s_in2(42,33),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(33)
		);
	s_in1(42,33)            <= s_out1(43,33);
	s_in2(42,33)            <= s_out2(43,34);
	s_locks_lower_in(42,33) <= s_locks_lower_out(43,33);

		normal_cell_42_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,34),
			fetch              => s_fetch(42,34),
			data_in            => s_data_in(42,34),
			data_out           => s_data_out(42,34),
			out1               => s_out1(42,34),
			out2               => s_out2(42,34),
			lock_lower_row_out => s_locks_lower_out(42,34),
			lock_lower_row_in  => s_locks_lower_in(42,34),
			in1                => s_in1(42,34),
			in2                => s_in2(42,34),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(34)
		);
	s_in1(42,34)            <= s_out1(43,34);
	s_in2(42,34)            <= s_out2(43,35);
	s_locks_lower_in(42,34) <= s_locks_lower_out(43,34);

		normal_cell_42_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,35),
			fetch              => s_fetch(42,35),
			data_in            => s_data_in(42,35),
			data_out           => s_data_out(42,35),
			out1               => s_out1(42,35),
			out2               => s_out2(42,35),
			lock_lower_row_out => s_locks_lower_out(42,35),
			lock_lower_row_in  => s_locks_lower_in(42,35),
			in1                => s_in1(42,35),
			in2                => s_in2(42,35),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(35)
		);
	s_in1(42,35)            <= s_out1(43,35);
	s_in2(42,35)            <= s_out2(43,36);
	s_locks_lower_in(42,35) <= s_locks_lower_out(43,35);

		normal_cell_42_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,36),
			fetch              => s_fetch(42,36),
			data_in            => s_data_in(42,36),
			data_out           => s_data_out(42,36),
			out1               => s_out1(42,36),
			out2               => s_out2(42,36),
			lock_lower_row_out => s_locks_lower_out(42,36),
			lock_lower_row_in  => s_locks_lower_in(42,36),
			in1                => s_in1(42,36),
			in2                => s_in2(42,36),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(36)
		);
	s_in1(42,36)            <= s_out1(43,36);
	s_in2(42,36)            <= s_out2(43,37);
	s_locks_lower_in(42,36) <= s_locks_lower_out(43,36);

		normal_cell_42_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,37),
			fetch              => s_fetch(42,37),
			data_in            => s_data_in(42,37),
			data_out           => s_data_out(42,37),
			out1               => s_out1(42,37),
			out2               => s_out2(42,37),
			lock_lower_row_out => s_locks_lower_out(42,37),
			lock_lower_row_in  => s_locks_lower_in(42,37),
			in1                => s_in1(42,37),
			in2                => s_in2(42,37),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(37)
		);
	s_in1(42,37)            <= s_out1(43,37);
	s_in2(42,37)            <= s_out2(43,38);
	s_locks_lower_in(42,37) <= s_locks_lower_out(43,37);

		normal_cell_42_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,38),
			fetch              => s_fetch(42,38),
			data_in            => s_data_in(42,38),
			data_out           => s_data_out(42,38),
			out1               => s_out1(42,38),
			out2               => s_out2(42,38),
			lock_lower_row_out => s_locks_lower_out(42,38),
			lock_lower_row_in  => s_locks_lower_in(42,38),
			in1                => s_in1(42,38),
			in2                => s_in2(42,38),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(38)
		);
	s_in1(42,38)            <= s_out1(43,38);
	s_in2(42,38)            <= s_out2(43,39);
	s_locks_lower_in(42,38) <= s_locks_lower_out(43,38);

		normal_cell_42_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,39),
			fetch              => s_fetch(42,39),
			data_in            => s_data_in(42,39),
			data_out           => s_data_out(42,39),
			out1               => s_out1(42,39),
			out2               => s_out2(42,39),
			lock_lower_row_out => s_locks_lower_out(42,39),
			lock_lower_row_in  => s_locks_lower_in(42,39),
			in1                => s_in1(42,39),
			in2                => s_in2(42,39),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(39)
		);
	s_in1(42,39)            <= s_out1(43,39);
	s_in2(42,39)            <= s_out2(43,40);
	s_locks_lower_in(42,39) <= s_locks_lower_out(43,39);

		normal_cell_42_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,40),
			fetch              => s_fetch(42,40),
			data_in            => s_data_in(42,40),
			data_out           => s_data_out(42,40),
			out1               => s_out1(42,40),
			out2               => s_out2(42,40),
			lock_lower_row_out => s_locks_lower_out(42,40),
			lock_lower_row_in  => s_locks_lower_in(42,40),
			in1                => s_in1(42,40),
			in2                => s_in2(42,40),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(40)
		);
	s_in1(42,40)            <= s_out1(43,40);
	s_in2(42,40)            <= s_out2(43,41);
	s_locks_lower_in(42,40) <= s_locks_lower_out(43,40);

		normal_cell_42_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,41),
			fetch              => s_fetch(42,41),
			data_in            => s_data_in(42,41),
			data_out           => s_data_out(42,41),
			out1               => s_out1(42,41),
			out2               => s_out2(42,41),
			lock_lower_row_out => s_locks_lower_out(42,41),
			lock_lower_row_in  => s_locks_lower_in(42,41),
			in1                => s_in1(42,41),
			in2                => s_in2(42,41),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(41)
		);
	s_in1(42,41)            <= s_out1(43,41);
	s_in2(42,41)            <= s_out2(43,42);
	s_locks_lower_in(42,41) <= s_locks_lower_out(43,41);

		normal_cell_42_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,42),
			fetch              => s_fetch(42,42),
			data_in            => s_data_in(42,42),
			data_out           => s_data_out(42,42),
			out1               => s_out1(42,42),
			out2               => s_out2(42,42),
			lock_lower_row_out => s_locks_lower_out(42,42),
			lock_lower_row_in  => s_locks_lower_in(42,42),
			in1                => s_in1(42,42),
			in2                => s_in2(42,42),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(42)
		);
	s_in1(42,42)            <= s_out1(43,42);
	s_in2(42,42)            <= s_out2(43,43);
	s_locks_lower_in(42,42) <= s_locks_lower_out(43,42);

		normal_cell_42_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,43),
			fetch              => s_fetch(42,43),
			data_in            => s_data_in(42,43),
			data_out           => s_data_out(42,43),
			out1               => s_out1(42,43),
			out2               => s_out2(42,43),
			lock_lower_row_out => s_locks_lower_out(42,43),
			lock_lower_row_in  => s_locks_lower_in(42,43),
			in1                => s_in1(42,43),
			in2                => s_in2(42,43),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(43)
		);
	s_in1(42,43)            <= s_out1(43,43);
	s_in2(42,43)            <= s_out2(43,44);
	s_locks_lower_in(42,43) <= s_locks_lower_out(43,43);

		normal_cell_42_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,44),
			fetch              => s_fetch(42,44),
			data_in            => s_data_in(42,44),
			data_out           => s_data_out(42,44),
			out1               => s_out1(42,44),
			out2               => s_out2(42,44),
			lock_lower_row_out => s_locks_lower_out(42,44),
			lock_lower_row_in  => s_locks_lower_in(42,44),
			in1                => s_in1(42,44),
			in2                => s_in2(42,44),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(44)
		);
	s_in1(42,44)            <= s_out1(43,44);
	s_in2(42,44)            <= s_out2(43,45);
	s_locks_lower_in(42,44) <= s_locks_lower_out(43,44);

		normal_cell_42_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,45),
			fetch              => s_fetch(42,45),
			data_in            => s_data_in(42,45),
			data_out           => s_data_out(42,45),
			out1               => s_out1(42,45),
			out2               => s_out2(42,45),
			lock_lower_row_out => s_locks_lower_out(42,45),
			lock_lower_row_in  => s_locks_lower_in(42,45),
			in1                => s_in1(42,45),
			in2                => s_in2(42,45),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(45)
		);
	s_in1(42,45)            <= s_out1(43,45);
	s_in2(42,45)            <= s_out2(43,46);
	s_locks_lower_in(42,45) <= s_locks_lower_out(43,45);

		normal_cell_42_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,46),
			fetch              => s_fetch(42,46),
			data_in            => s_data_in(42,46),
			data_out           => s_data_out(42,46),
			out1               => s_out1(42,46),
			out2               => s_out2(42,46),
			lock_lower_row_out => s_locks_lower_out(42,46),
			lock_lower_row_in  => s_locks_lower_in(42,46),
			in1                => s_in1(42,46),
			in2                => s_in2(42,46),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(46)
		);
	s_in1(42,46)            <= s_out1(43,46);
	s_in2(42,46)            <= s_out2(43,47);
	s_locks_lower_in(42,46) <= s_locks_lower_out(43,46);

		normal_cell_42_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,47),
			fetch              => s_fetch(42,47),
			data_in            => s_data_in(42,47),
			data_out           => s_data_out(42,47),
			out1               => s_out1(42,47),
			out2               => s_out2(42,47),
			lock_lower_row_out => s_locks_lower_out(42,47),
			lock_lower_row_in  => s_locks_lower_in(42,47),
			in1                => s_in1(42,47),
			in2                => s_in2(42,47),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(47)
		);
	s_in1(42,47)            <= s_out1(43,47);
	s_in2(42,47)            <= s_out2(43,48);
	s_locks_lower_in(42,47) <= s_locks_lower_out(43,47);

		normal_cell_42_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,48),
			fetch              => s_fetch(42,48),
			data_in            => s_data_in(42,48),
			data_out           => s_data_out(42,48),
			out1               => s_out1(42,48),
			out2               => s_out2(42,48),
			lock_lower_row_out => s_locks_lower_out(42,48),
			lock_lower_row_in  => s_locks_lower_in(42,48),
			in1                => s_in1(42,48),
			in2                => s_in2(42,48),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(48)
		);
	s_in1(42,48)            <= s_out1(43,48);
	s_in2(42,48)            <= s_out2(43,49);
	s_locks_lower_in(42,48) <= s_locks_lower_out(43,48);

		normal_cell_42_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,49),
			fetch              => s_fetch(42,49),
			data_in            => s_data_in(42,49),
			data_out           => s_data_out(42,49),
			out1               => s_out1(42,49),
			out2               => s_out2(42,49),
			lock_lower_row_out => s_locks_lower_out(42,49),
			lock_lower_row_in  => s_locks_lower_in(42,49),
			in1                => s_in1(42,49),
			in2                => s_in2(42,49),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(49)
		);
	s_in1(42,49)            <= s_out1(43,49);
	s_in2(42,49)            <= s_out2(43,50);
	s_locks_lower_in(42,49) <= s_locks_lower_out(43,49);

		normal_cell_42_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,50),
			fetch              => s_fetch(42,50),
			data_in            => s_data_in(42,50),
			data_out           => s_data_out(42,50),
			out1               => s_out1(42,50),
			out2               => s_out2(42,50),
			lock_lower_row_out => s_locks_lower_out(42,50),
			lock_lower_row_in  => s_locks_lower_in(42,50),
			in1                => s_in1(42,50),
			in2                => s_in2(42,50),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(50)
		);
	s_in1(42,50)            <= s_out1(43,50);
	s_in2(42,50)            <= s_out2(43,51);
	s_locks_lower_in(42,50) <= s_locks_lower_out(43,50);

		normal_cell_42_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,51),
			fetch              => s_fetch(42,51),
			data_in            => s_data_in(42,51),
			data_out           => s_data_out(42,51),
			out1               => s_out1(42,51),
			out2               => s_out2(42,51),
			lock_lower_row_out => s_locks_lower_out(42,51),
			lock_lower_row_in  => s_locks_lower_in(42,51),
			in1                => s_in1(42,51),
			in2                => s_in2(42,51),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(51)
		);
	s_in1(42,51)            <= s_out1(43,51);
	s_in2(42,51)            <= s_out2(43,52);
	s_locks_lower_in(42,51) <= s_locks_lower_out(43,51);

		normal_cell_42_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,52),
			fetch              => s_fetch(42,52),
			data_in            => s_data_in(42,52),
			data_out           => s_data_out(42,52),
			out1               => s_out1(42,52),
			out2               => s_out2(42,52),
			lock_lower_row_out => s_locks_lower_out(42,52),
			lock_lower_row_in  => s_locks_lower_in(42,52),
			in1                => s_in1(42,52),
			in2                => s_in2(42,52),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(52)
		);
	s_in1(42,52)            <= s_out1(43,52);
	s_in2(42,52)            <= s_out2(43,53);
	s_locks_lower_in(42,52) <= s_locks_lower_out(43,52);

		normal_cell_42_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,53),
			fetch              => s_fetch(42,53),
			data_in            => s_data_in(42,53),
			data_out           => s_data_out(42,53),
			out1               => s_out1(42,53),
			out2               => s_out2(42,53),
			lock_lower_row_out => s_locks_lower_out(42,53),
			lock_lower_row_in  => s_locks_lower_in(42,53),
			in1                => s_in1(42,53),
			in2                => s_in2(42,53),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(53)
		);
	s_in1(42,53)            <= s_out1(43,53);
	s_in2(42,53)            <= s_out2(43,54);
	s_locks_lower_in(42,53) <= s_locks_lower_out(43,53);

		normal_cell_42_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,54),
			fetch              => s_fetch(42,54),
			data_in            => s_data_in(42,54),
			data_out           => s_data_out(42,54),
			out1               => s_out1(42,54),
			out2               => s_out2(42,54),
			lock_lower_row_out => s_locks_lower_out(42,54),
			lock_lower_row_in  => s_locks_lower_in(42,54),
			in1                => s_in1(42,54),
			in2                => s_in2(42,54),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(54)
		);
	s_in1(42,54)            <= s_out1(43,54);
	s_in2(42,54)            <= s_out2(43,55);
	s_locks_lower_in(42,54) <= s_locks_lower_out(43,54);

		normal_cell_42_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,55),
			fetch              => s_fetch(42,55),
			data_in            => s_data_in(42,55),
			data_out           => s_data_out(42,55),
			out1               => s_out1(42,55),
			out2               => s_out2(42,55),
			lock_lower_row_out => s_locks_lower_out(42,55),
			lock_lower_row_in  => s_locks_lower_in(42,55),
			in1                => s_in1(42,55),
			in2                => s_in2(42,55),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(55)
		);
	s_in1(42,55)            <= s_out1(43,55);
	s_in2(42,55)            <= s_out2(43,56);
	s_locks_lower_in(42,55) <= s_locks_lower_out(43,55);

		normal_cell_42_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,56),
			fetch              => s_fetch(42,56),
			data_in            => s_data_in(42,56),
			data_out           => s_data_out(42,56),
			out1               => s_out1(42,56),
			out2               => s_out2(42,56),
			lock_lower_row_out => s_locks_lower_out(42,56),
			lock_lower_row_in  => s_locks_lower_in(42,56),
			in1                => s_in1(42,56),
			in2                => s_in2(42,56),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(56)
		);
	s_in1(42,56)            <= s_out1(43,56);
	s_in2(42,56)            <= s_out2(43,57);
	s_locks_lower_in(42,56) <= s_locks_lower_out(43,56);

		normal_cell_42_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,57),
			fetch              => s_fetch(42,57),
			data_in            => s_data_in(42,57),
			data_out           => s_data_out(42,57),
			out1               => s_out1(42,57),
			out2               => s_out2(42,57),
			lock_lower_row_out => s_locks_lower_out(42,57),
			lock_lower_row_in  => s_locks_lower_in(42,57),
			in1                => s_in1(42,57),
			in2                => s_in2(42,57),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(57)
		);
	s_in1(42,57)            <= s_out1(43,57);
	s_in2(42,57)            <= s_out2(43,58);
	s_locks_lower_in(42,57) <= s_locks_lower_out(43,57);

		normal_cell_42_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,58),
			fetch              => s_fetch(42,58),
			data_in            => s_data_in(42,58),
			data_out           => s_data_out(42,58),
			out1               => s_out1(42,58),
			out2               => s_out2(42,58),
			lock_lower_row_out => s_locks_lower_out(42,58),
			lock_lower_row_in  => s_locks_lower_in(42,58),
			in1                => s_in1(42,58),
			in2                => s_in2(42,58),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(58)
		);
	s_in1(42,58)            <= s_out1(43,58);
	s_in2(42,58)            <= s_out2(43,59);
	s_locks_lower_in(42,58) <= s_locks_lower_out(43,58);

		normal_cell_42_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,59),
			fetch              => s_fetch(42,59),
			data_in            => s_data_in(42,59),
			data_out           => s_data_out(42,59),
			out1               => s_out1(42,59),
			out2               => s_out2(42,59),
			lock_lower_row_out => s_locks_lower_out(42,59),
			lock_lower_row_in  => s_locks_lower_in(42,59),
			in1                => s_in1(42,59),
			in2                => s_in2(42,59),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(59)
		);
	s_in1(42,59)            <= s_out1(43,59);
	s_in2(42,59)            <= s_out2(43,60);
	s_locks_lower_in(42,59) <= s_locks_lower_out(43,59);

		last_col_cell_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(42,60),
			fetch              => s_fetch(42,60),
			data_in            => s_data_in(42,60),
			data_out           => s_data_out(42,60),
			out1               => s_out1(42,60),
			out2               => s_out2(42,60),
			lock_lower_row_out => s_locks_lower_out(42,60),
			lock_lower_row_in  => s_locks_lower_in(42,60),
			in1                => s_in1(42,60),
			in2                => (others => '0'),
			lock_row           => s_locks(42),
			piv_found          => s_piv_found,
			row_data           => s_row_data(42),
			col_data           => s_col_data(60)
		);
	s_in1(42,60)            <= s_out1(43,60);
	s_locks_lower_in(42,60) <= s_locks_lower_out(43,60);

		normal_cell_43_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,1),
			fetch              => s_fetch(43,1),
			data_in            => s_data_in(43,1),
			data_out           => s_data_out(43,1),
			out1               => s_out1(43,1),
			out2               => s_out2(43,1),
			lock_lower_row_out => s_locks_lower_out(43,1),
			lock_lower_row_in  => s_locks_lower_in(43,1),
			in1                => s_in1(43,1),
			in2                => s_in2(43,1),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(1)
		);
	s_in1(43,1)            <= s_out1(44,1);
	s_in2(43,1)            <= s_out2(44,2);
	s_locks_lower_in(43,1) <= s_locks_lower_out(44,1);

		normal_cell_43_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,2),
			fetch              => s_fetch(43,2),
			data_in            => s_data_in(43,2),
			data_out           => s_data_out(43,2),
			out1               => s_out1(43,2),
			out2               => s_out2(43,2),
			lock_lower_row_out => s_locks_lower_out(43,2),
			lock_lower_row_in  => s_locks_lower_in(43,2),
			in1                => s_in1(43,2),
			in2                => s_in2(43,2),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(2)
		);
	s_in1(43,2)            <= s_out1(44,2);
	s_in2(43,2)            <= s_out2(44,3);
	s_locks_lower_in(43,2) <= s_locks_lower_out(44,2);

		normal_cell_43_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,3),
			fetch              => s_fetch(43,3),
			data_in            => s_data_in(43,3),
			data_out           => s_data_out(43,3),
			out1               => s_out1(43,3),
			out2               => s_out2(43,3),
			lock_lower_row_out => s_locks_lower_out(43,3),
			lock_lower_row_in  => s_locks_lower_in(43,3),
			in1                => s_in1(43,3),
			in2                => s_in2(43,3),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(3)
		);
	s_in1(43,3)            <= s_out1(44,3);
	s_in2(43,3)            <= s_out2(44,4);
	s_locks_lower_in(43,3) <= s_locks_lower_out(44,3);

		normal_cell_43_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,4),
			fetch              => s_fetch(43,4),
			data_in            => s_data_in(43,4),
			data_out           => s_data_out(43,4),
			out1               => s_out1(43,4),
			out2               => s_out2(43,4),
			lock_lower_row_out => s_locks_lower_out(43,4),
			lock_lower_row_in  => s_locks_lower_in(43,4),
			in1                => s_in1(43,4),
			in2                => s_in2(43,4),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(4)
		);
	s_in1(43,4)            <= s_out1(44,4);
	s_in2(43,4)            <= s_out2(44,5);
	s_locks_lower_in(43,4) <= s_locks_lower_out(44,4);

		normal_cell_43_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,5),
			fetch              => s_fetch(43,5),
			data_in            => s_data_in(43,5),
			data_out           => s_data_out(43,5),
			out1               => s_out1(43,5),
			out2               => s_out2(43,5),
			lock_lower_row_out => s_locks_lower_out(43,5),
			lock_lower_row_in  => s_locks_lower_in(43,5),
			in1                => s_in1(43,5),
			in2                => s_in2(43,5),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(5)
		);
	s_in1(43,5)            <= s_out1(44,5);
	s_in2(43,5)            <= s_out2(44,6);
	s_locks_lower_in(43,5) <= s_locks_lower_out(44,5);

		normal_cell_43_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,6),
			fetch              => s_fetch(43,6),
			data_in            => s_data_in(43,6),
			data_out           => s_data_out(43,6),
			out1               => s_out1(43,6),
			out2               => s_out2(43,6),
			lock_lower_row_out => s_locks_lower_out(43,6),
			lock_lower_row_in  => s_locks_lower_in(43,6),
			in1                => s_in1(43,6),
			in2                => s_in2(43,6),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(6)
		);
	s_in1(43,6)            <= s_out1(44,6);
	s_in2(43,6)            <= s_out2(44,7);
	s_locks_lower_in(43,6) <= s_locks_lower_out(44,6);

		normal_cell_43_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,7),
			fetch              => s_fetch(43,7),
			data_in            => s_data_in(43,7),
			data_out           => s_data_out(43,7),
			out1               => s_out1(43,7),
			out2               => s_out2(43,7),
			lock_lower_row_out => s_locks_lower_out(43,7),
			lock_lower_row_in  => s_locks_lower_in(43,7),
			in1                => s_in1(43,7),
			in2                => s_in2(43,7),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(7)
		);
	s_in1(43,7)            <= s_out1(44,7);
	s_in2(43,7)            <= s_out2(44,8);
	s_locks_lower_in(43,7) <= s_locks_lower_out(44,7);

		normal_cell_43_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,8),
			fetch              => s_fetch(43,8),
			data_in            => s_data_in(43,8),
			data_out           => s_data_out(43,8),
			out1               => s_out1(43,8),
			out2               => s_out2(43,8),
			lock_lower_row_out => s_locks_lower_out(43,8),
			lock_lower_row_in  => s_locks_lower_in(43,8),
			in1                => s_in1(43,8),
			in2                => s_in2(43,8),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(8)
		);
	s_in1(43,8)            <= s_out1(44,8);
	s_in2(43,8)            <= s_out2(44,9);
	s_locks_lower_in(43,8) <= s_locks_lower_out(44,8);

		normal_cell_43_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,9),
			fetch              => s_fetch(43,9),
			data_in            => s_data_in(43,9),
			data_out           => s_data_out(43,9),
			out1               => s_out1(43,9),
			out2               => s_out2(43,9),
			lock_lower_row_out => s_locks_lower_out(43,9),
			lock_lower_row_in  => s_locks_lower_in(43,9),
			in1                => s_in1(43,9),
			in2                => s_in2(43,9),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(9)
		);
	s_in1(43,9)            <= s_out1(44,9);
	s_in2(43,9)            <= s_out2(44,10);
	s_locks_lower_in(43,9) <= s_locks_lower_out(44,9);

		normal_cell_43_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,10),
			fetch              => s_fetch(43,10),
			data_in            => s_data_in(43,10),
			data_out           => s_data_out(43,10),
			out1               => s_out1(43,10),
			out2               => s_out2(43,10),
			lock_lower_row_out => s_locks_lower_out(43,10),
			lock_lower_row_in  => s_locks_lower_in(43,10),
			in1                => s_in1(43,10),
			in2                => s_in2(43,10),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(10)
		);
	s_in1(43,10)            <= s_out1(44,10);
	s_in2(43,10)            <= s_out2(44,11);
	s_locks_lower_in(43,10) <= s_locks_lower_out(44,10);

		normal_cell_43_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,11),
			fetch              => s_fetch(43,11),
			data_in            => s_data_in(43,11),
			data_out           => s_data_out(43,11),
			out1               => s_out1(43,11),
			out2               => s_out2(43,11),
			lock_lower_row_out => s_locks_lower_out(43,11),
			lock_lower_row_in  => s_locks_lower_in(43,11),
			in1                => s_in1(43,11),
			in2                => s_in2(43,11),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(11)
		);
	s_in1(43,11)            <= s_out1(44,11);
	s_in2(43,11)            <= s_out2(44,12);
	s_locks_lower_in(43,11) <= s_locks_lower_out(44,11);

		normal_cell_43_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,12),
			fetch              => s_fetch(43,12),
			data_in            => s_data_in(43,12),
			data_out           => s_data_out(43,12),
			out1               => s_out1(43,12),
			out2               => s_out2(43,12),
			lock_lower_row_out => s_locks_lower_out(43,12),
			lock_lower_row_in  => s_locks_lower_in(43,12),
			in1                => s_in1(43,12),
			in2                => s_in2(43,12),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(12)
		);
	s_in1(43,12)            <= s_out1(44,12);
	s_in2(43,12)            <= s_out2(44,13);
	s_locks_lower_in(43,12) <= s_locks_lower_out(44,12);

		normal_cell_43_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,13),
			fetch              => s_fetch(43,13),
			data_in            => s_data_in(43,13),
			data_out           => s_data_out(43,13),
			out1               => s_out1(43,13),
			out2               => s_out2(43,13),
			lock_lower_row_out => s_locks_lower_out(43,13),
			lock_lower_row_in  => s_locks_lower_in(43,13),
			in1                => s_in1(43,13),
			in2                => s_in2(43,13),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(13)
		);
	s_in1(43,13)            <= s_out1(44,13);
	s_in2(43,13)            <= s_out2(44,14);
	s_locks_lower_in(43,13) <= s_locks_lower_out(44,13);

		normal_cell_43_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,14),
			fetch              => s_fetch(43,14),
			data_in            => s_data_in(43,14),
			data_out           => s_data_out(43,14),
			out1               => s_out1(43,14),
			out2               => s_out2(43,14),
			lock_lower_row_out => s_locks_lower_out(43,14),
			lock_lower_row_in  => s_locks_lower_in(43,14),
			in1                => s_in1(43,14),
			in2                => s_in2(43,14),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(14)
		);
	s_in1(43,14)            <= s_out1(44,14);
	s_in2(43,14)            <= s_out2(44,15);
	s_locks_lower_in(43,14) <= s_locks_lower_out(44,14);

		normal_cell_43_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,15),
			fetch              => s_fetch(43,15),
			data_in            => s_data_in(43,15),
			data_out           => s_data_out(43,15),
			out1               => s_out1(43,15),
			out2               => s_out2(43,15),
			lock_lower_row_out => s_locks_lower_out(43,15),
			lock_lower_row_in  => s_locks_lower_in(43,15),
			in1                => s_in1(43,15),
			in2                => s_in2(43,15),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(15)
		);
	s_in1(43,15)            <= s_out1(44,15);
	s_in2(43,15)            <= s_out2(44,16);
	s_locks_lower_in(43,15) <= s_locks_lower_out(44,15);

		normal_cell_43_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,16),
			fetch              => s_fetch(43,16),
			data_in            => s_data_in(43,16),
			data_out           => s_data_out(43,16),
			out1               => s_out1(43,16),
			out2               => s_out2(43,16),
			lock_lower_row_out => s_locks_lower_out(43,16),
			lock_lower_row_in  => s_locks_lower_in(43,16),
			in1                => s_in1(43,16),
			in2                => s_in2(43,16),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(16)
		);
	s_in1(43,16)            <= s_out1(44,16);
	s_in2(43,16)            <= s_out2(44,17);
	s_locks_lower_in(43,16) <= s_locks_lower_out(44,16);

		normal_cell_43_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,17),
			fetch              => s_fetch(43,17),
			data_in            => s_data_in(43,17),
			data_out           => s_data_out(43,17),
			out1               => s_out1(43,17),
			out2               => s_out2(43,17),
			lock_lower_row_out => s_locks_lower_out(43,17),
			lock_lower_row_in  => s_locks_lower_in(43,17),
			in1                => s_in1(43,17),
			in2                => s_in2(43,17),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(17)
		);
	s_in1(43,17)            <= s_out1(44,17);
	s_in2(43,17)            <= s_out2(44,18);
	s_locks_lower_in(43,17) <= s_locks_lower_out(44,17);

		normal_cell_43_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,18),
			fetch              => s_fetch(43,18),
			data_in            => s_data_in(43,18),
			data_out           => s_data_out(43,18),
			out1               => s_out1(43,18),
			out2               => s_out2(43,18),
			lock_lower_row_out => s_locks_lower_out(43,18),
			lock_lower_row_in  => s_locks_lower_in(43,18),
			in1                => s_in1(43,18),
			in2                => s_in2(43,18),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(18)
		);
	s_in1(43,18)            <= s_out1(44,18);
	s_in2(43,18)            <= s_out2(44,19);
	s_locks_lower_in(43,18) <= s_locks_lower_out(44,18);

		normal_cell_43_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,19),
			fetch              => s_fetch(43,19),
			data_in            => s_data_in(43,19),
			data_out           => s_data_out(43,19),
			out1               => s_out1(43,19),
			out2               => s_out2(43,19),
			lock_lower_row_out => s_locks_lower_out(43,19),
			lock_lower_row_in  => s_locks_lower_in(43,19),
			in1                => s_in1(43,19),
			in2                => s_in2(43,19),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(19)
		);
	s_in1(43,19)            <= s_out1(44,19);
	s_in2(43,19)            <= s_out2(44,20);
	s_locks_lower_in(43,19) <= s_locks_lower_out(44,19);

		normal_cell_43_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,20),
			fetch              => s_fetch(43,20),
			data_in            => s_data_in(43,20),
			data_out           => s_data_out(43,20),
			out1               => s_out1(43,20),
			out2               => s_out2(43,20),
			lock_lower_row_out => s_locks_lower_out(43,20),
			lock_lower_row_in  => s_locks_lower_in(43,20),
			in1                => s_in1(43,20),
			in2                => s_in2(43,20),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(20)
		);
	s_in1(43,20)            <= s_out1(44,20);
	s_in2(43,20)            <= s_out2(44,21);
	s_locks_lower_in(43,20) <= s_locks_lower_out(44,20);

		normal_cell_43_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,21),
			fetch              => s_fetch(43,21),
			data_in            => s_data_in(43,21),
			data_out           => s_data_out(43,21),
			out1               => s_out1(43,21),
			out2               => s_out2(43,21),
			lock_lower_row_out => s_locks_lower_out(43,21),
			lock_lower_row_in  => s_locks_lower_in(43,21),
			in1                => s_in1(43,21),
			in2                => s_in2(43,21),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(21)
		);
	s_in1(43,21)            <= s_out1(44,21);
	s_in2(43,21)            <= s_out2(44,22);
	s_locks_lower_in(43,21) <= s_locks_lower_out(44,21);

		normal_cell_43_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,22),
			fetch              => s_fetch(43,22),
			data_in            => s_data_in(43,22),
			data_out           => s_data_out(43,22),
			out1               => s_out1(43,22),
			out2               => s_out2(43,22),
			lock_lower_row_out => s_locks_lower_out(43,22),
			lock_lower_row_in  => s_locks_lower_in(43,22),
			in1                => s_in1(43,22),
			in2                => s_in2(43,22),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(22)
		);
	s_in1(43,22)            <= s_out1(44,22);
	s_in2(43,22)            <= s_out2(44,23);
	s_locks_lower_in(43,22) <= s_locks_lower_out(44,22);

		normal_cell_43_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,23),
			fetch              => s_fetch(43,23),
			data_in            => s_data_in(43,23),
			data_out           => s_data_out(43,23),
			out1               => s_out1(43,23),
			out2               => s_out2(43,23),
			lock_lower_row_out => s_locks_lower_out(43,23),
			lock_lower_row_in  => s_locks_lower_in(43,23),
			in1                => s_in1(43,23),
			in2                => s_in2(43,23),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(23)
		);
	s_in1(43,23)            <= s_out1(44,23);
	s_in2(43,23)            <= s_out2(44,24);
	s_locks_lower_in(43,23) <= s_locks_lower_out(44,23);

		normal_cell_43_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,24),
			fetch              => s_fetch(43,24),
			data_in            => s_data_in(43,24),
			data_out           => s_data_out(43,24),
			out1               => s_out1(43,24),
			out2               => s_out2(43,24),
			lock_lower_row_out => s_locks_lower_out(43,24),
			lock_lower_row_in  => s_locks_lower_in(43,24),
			in1                => s_in1(43,24),
			in2                => s_in2(43,24),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(24)
		);
	s_in1(43,24)            <= s_out1(44,24);
	s_in2(43,24)            <= s_out2(44,25);
	s_locks_lower_in(43,24) <= s_locks_lower_out(44,24);

		normal_cell_43_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,25),
			fetch              => s_fetch(43,25),
			data_in            => s_data_in(43,25),
			data_out           => s_data_out(43,25),
			out1               => s_out1(43,25),
			out2               => s_out2(43,25),
			lock_lower_row_out => s_locks_lower_out(43,25),
			lock_lower_row_in  => s_locks_lower_in(43,25),
			in1                => s_in1(43,25),
			in2                => s_in2(43,25),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(25)
		);
	s_in1(43,25)            <= s_out1(44,25);
	s_in2(43,25)            <= s_out2(44,26);
	s_locks_lower_in(43,25) <= s_locks_lower_out(44,25);

		normal_cell_43_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,26),
			fetch              => s_fetch(43,26),
			data_in            => s_data_in(43,26),
			data_out           => s_data_out(43,26),
			out1               => s_out1(43,26),
			out2               => s_out2(43,26),
			lock_lower_row_out => s_locks_lower_out(43,26),
			lock_lower_row_in  => s_locks_lower_in(43,26),
			in1                => s_in1(43,26),
			in2                => s_in2(43,26),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(26)
		);
	s_in1(43,26)            <= s_out1(44,26);
	s_in2(43,26)            <= s_out2(44,27);
	s_locks_lower_in(43,26) <= s_locks_lower_out(44,26);

		normal_cell_43_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,27),
			fetch              => s_fetch(43,27),
			data_in            => s_data_in(43,27),
			data_out           => s_data_out(43,27),
			out1               => s_out1(43,27),
			out2               => s_out2(43,27),
			lock_lower_row_out => s_locks_lower_out(43,27),
			lock_lower_row_in  => s_locks_lower_in(43,27),
			in1                => s_in1(43,27),
			in2                => s_in2(43,27),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(27)
		);
	s_in1(43,27)            <= s_out1(44,27);
	s_in2(43,27)            <= s_out2(44,28);
	s_locks_lower_in(43,27) <= s_locks_lower_out(44,27);

		normal_cell_43_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,28),
			fetch              => s_fetch(43,28),
			data_in            => s_data_in(43,28),
			data_out           => s_data_out(43,28),
			out1               => s_out1(43,28),
			out2               => s_out2(43,28),
			lock_lower_row_out => s_locks_lower_out(43,28),
			lock_lower_row_in  => s_locks_lower_in(43,28),
			in1                => s_in1(43,28),
			in2                => s_in2(43,28),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(28)
		);
	s_in1(43,28)            <= s_out1(44,28);
	s_in2(43,28)            <= s_out2(44,29);
	s_locks_lower_in(43,28) <= s_locks_lower_out(44,28);

		normal_cell_43_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,29),
			fetch              => s_fetch(43,29),
			data_in            => s_data_in(43,29),
			data_out           => s_data_out(43,29),
			out1               => s_out1(43,29),
			out2               => s_out2(43,29),
			lock_lower_row_out => s_locks_lower_out(43,29),
			lock_lower_row_in  => s_locks_lower_in(43,29),
			in1                => s_in1(43,29),
			in2                => s_in2(43,29),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(29)
		);
	s_in1(43,29)            <= s_out1(44,29);
	s_in2(43,29)            <= s_out2(44,30);
	s_locks_lower_in(43,29) <= s_locks_lower_out(44,29);

		normal_cell_43_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,30),
			fetch              => s_fetch(43,30),
			data_in            => s_data_in(43,30),
			data_out           => s_data_out(43,30),
			out1               => s_out1(43,30),
			out2               => s_out2(43,30),
			lock_lower_row_out => s_locks_lower_out(43,30),
			lock_lower_row_in  => s_locks_lower_in(43,30),
			in1                => s_in1(43,30),
			in2                => s_in2(43,30),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(30)
		);
	s_in1(43,30)            <= s_out1(44,30);
	s_in2(43,30)            <= s_out2(44,31);
	s_locks_lower_in(43,30) <= s_locks_lower_out(44,30);

		normal_cell_43_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,31),
			fetch              => s_fetch(43,31),
			data_in            => s_data_in(43,31),
			data_out           => s_data_out(43,31),
			out1               => s_out1(43,31),
			out2               => s_out2(43,31),
			lock_lower_row_out => s_locks_lower_out(43,31),
			lock_lower_row_in  => s_locks_lower_in(43,31),
			in1                => s_in1(43,31),
			in2                => s_in2(43,31),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(31)
		);
	s_in1(43,31)            <= s_out1(44,31);
	s_in2(43,31)            <= s_out2(44,32);
	s_locks_lower_in(43,31) <= s_locks_lower_out(44,31);

		normal_cell_43_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,32),
			fetch              => s_fetch(43,32),
			data_in            => s_data_in(43,32),
			data_out           => s_data_out(43,32),
			out1               => s_out1(43,32),
			out2               => s_out2(43,32),
			lock_lower_row_out => s_locks_lower_out(43,32),
			lock_lower_row_in  => s_locks_lower_in(43,32),
			in1                => s_in1(43,32),
			in2                => s_in2(43,32),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(32)
		);
	s_in1(43,32)            <= s_out1(44,32);
	s_in2(43,32)            <= s_out2(44,33);
	s_locks_lower_in(43,32) <= s_locks_lower_out(44,32);

		normal_cell_43_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,33),
			fetch              => s_fetch(43,33),
			data_in            => s_data_in(43,33),
			data_out           => s_data_out(43,33),
			out1               => s_out1(43,33),
			out2               => s_out2(43,33),
			lock_lower_row_out => s_locks_lower_out(43,33),
			lock_lower_row_in  => s_locks_lower_in(43,33),
			in1                => s_in1(43,33),
			in2                => s_in2(43,33),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(33)
		);
	s_in1(43,33)            <= s_out1(44,33);
	s_in2(43,33)            <= s_out2(44,34);
	s_locks_lower_in(43,33) <= s_locks_lower_out(44,33);

		normal_cell_43_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,34),
			fetch              => s_fetch(43,34),
			data_in            => s_data_in(43,34),
			data_out           => s_data_out(43,34),
			out1               => s_out1(43,34),
			out2               => s_out2(43,34),
			lock_lower_row_out => s_locks_lower_out(43,34),
			lock_lower_row_in  => s_locks_lower_in(43,34),
			in1                => s_in1(43,34),
			in2                => s_in2(43,34),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(34)
		);
	s_in1(43,34)            <= s_out1(44,34);
	s_in2(43,34)            <= s_out2(44,35);
	s_locks_lower_in(43,34) <= s_locks_lower_out(44,34);

		normal_cell_43_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,35),
			fetch              => s_fetch(43,35),
			data_in            => s_data_in(43,35),
			data_out           => s_data_out(43,35),
			out1               => s_out1(43,35),
			out2               => s_out2(43,35),
			lock_lower_row_out => s_locks_lower_out(43,35),
			lock_lower_row_in  => s_locks_lower_in(43,35),
			in1                => s_in1(43,35),
			in2                => s_in2(43,35),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(35)
		);
	s_in1(43,35)            <= s_out1(44,35);
	s_in2(43,35)            <= s_out2(44,36);
	s_locks_lower_in(43,35) <= s_locks_lower_out(44,35);

		normal_cell_43_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,36),
			fetch              => s_fetch(43,36),
			data_in            => s_data_in(43,36),
			data_out           => s_data_out(43,36),
			out1               => s_out1(43,36),
			out2               => s_out2(43,36),
			lock_lower_row_out => s_locks_lower_out(43,36),
			lock_lower_row_in  => s_locks_lower_in(43,36),
			in1                => s_in1(43,36),
			in2                => s_in2(43,36),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(36)
		);
	s_in1(43,36)            <= s_out1(44,36);
	s_in2(43,36)            <= s_out2(44,37);
	s_locks_lower_in(43,36) <= s_locks_lower_out(44,36);

		normal_cell_43_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,37),
			fetch              => s_fetch(43,37),
			data_in            => s_data_in(43,37),
			data_out           => s_data_out(43,37),
			out1               => s_out1(43,37),
			out2               => s_out2(43,37),
			lock_lower_row_out => s_locks_lower_out(43,37),
			lock_lower_row_in  => s_locks_lower_in(43,37),
			in1                => s_in1(43,37),
			in2                => s_in2(43,37),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(37)
		);
	s_in1(43,37)            <= s_out1(44,37);
	s_in2(43,37)            <= s_out2(44,38);
	s_locks_lower_in(43,37) <= s_locks_lower_out(44,37);

		normal_cell_43_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,38),
			fetch              => s_fetch(43,38),
			data_in            => s_data_in(43,38),
			data_out           => s_data_out(43,38),
			out1               => s_out1(43,38),
			out2               => s_out2(43,38),
			lock_lower_row_out => s_locks_lower_out(43,38),
			lock_lower_row_in  => s_locks_lower_in(43,38),
			in1                => s_in1(43,38),
			in2                => s_in2(43,38),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(38)
		);
	s_in1(43,38)            <= s_out1(44,38);
	s_in2(43,38)            <= s_out2(44,39);
	s_locks_lower_in(43,38) <= s_locks_lower_out(44,38);

		normal_cell_43_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,39),
			fetch              => s_fetch(43,39),
			data_in            => s_data_in(43,39),
			data_out           => s_data_out(43,39),
			out1               => s_out1(43,39),
			out2               => s_out2(43,39),
			lock_lower_row_out => s_locks_lower_out(43,39),
			lock_lower_row_in  => s_locks_lower_in(43,39),
			in1                => s_in1(43,39),
			in2                => s_in2(43,39),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(39)
		);
	s_in1(43,39)            <= s_out1(44,39);
	s_in2(43,39)            <= s_out2(44,40);
	s_locks_lower_in(43,39) <= s_locks_lower_out(44,39);

		normal_cell_43_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,40),
			fetch              => s_fetch(43,40),
			data_in            => s_data_in(43,40),
			data_out           => s_data_out(43,40),
			out1               => s_out1(43,40),
			out2               => s_out2(43,40),
			lock_lower_row_out => s_locks_lower_out(43,40),
			lock_lower_row_in  => s_locks_lower_in(43,40),
			in1                => s_in1(43,40),
			in2                => s_in2(43,40),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(40)
		);
	s_in1(43,40)            <= s_out1(44,40);
	s_in2(43,40)            <= s_out2(44,41);
	s_locks_lower_in(43,40) <= s_locks_lower_out(44,40);

		normal_cell_43_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,41),
			fetch              => s_fetch(43,41),
			data_in            => s_data_in(43,41),
			data_out           => s_data_out(43,41),
			out1               => s_out1(43,41),
			out2               => s_out2(43,41),
			lock_lower_row_out => s_locks_lower_out(43,41),
			lock_lower_row_in  => s_locks_lower_in(43,41),
			in1                => s_in1(43,41),
			in2                => s_in2(43,41),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(41)
		);
	s_in1(43,41)            <= s_out1(44,41);
	s_in2(43,41)            <= s_out2(44,42);
	s_locks_lower_in(43,41) <= s_locks_lower_out(44,41);

		normal_cell_43_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,42),
			fetch              => s_fetch(43,42),
			data_in            => s_data_in(43,42),
			data_out           => s_data_out(43,42),
			out1               => s_out1(43,42),
			out2               => s_out2(43,42),
			lock_lower_row_out => s_locks_lower_out(43,42),
			lock_lower_row_in  => s_locks_lower_in(43,42),
			in1                => s_in1(43,42),
			in2                => s_in2(43,42),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(42)
		);
	s_in1(43,42)            <= s_out1(44,42);
	s_in2(43,42)            <= s_out2(44,43);
	s_locks_lower_in(43,42) <= s_locks_lower_out(44,42);

		normal_cell_43_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,43),
			fetch              => s_fetch(43,43),
			data_in            => s_data_in(43,43),
			data_out           => s_data_out(43,43),
			out1               => s_out1(43,43),
			out2               => s_out2(43,43),
			lock_lower_row_out => s_locks_lower_out(43,43),
			lock_lower_row_in  => s_locks_lower_in(43,43),
			in1                => s_in1(43,43),
			in2                => s_in2(43,43),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(43)
		);
	s_in1(43,43)            <= s_out1(44,43);
	s_in2(43,43)            <= s_out2(44,44);
	s_locks_lower_in(43,43) <= s_locks_lower_out(44,43);

		normal_cell_43_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,44),
			fetch              => s_fetch(43,44),
			data_in            => s_data_in(43,44),
			data_out           => s_data_out(43,44),
			out1               => s_out1(43,44),
			out2               => s_out2(43,44),
			lock_lower_row_out => s_locks_lower_out(43,44),
			lock_lower_row_in  => s_locks_lower_in(43,44),
			in1                => s_in1(43,44),
			in2                => s_in2(43,44),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(44)
		);
	s_in1(43,44)            <= s_out1(44,44);
	s_in2(43,44)            <= s_out2(44,45);
	s_locks_lower_in(43,44) <= s_locks_lower_out(44,44);

		normal_cell_43_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,45),
			fetch              => s_fetch(43,45),
			data_in            => s_data_in(43,45),
			data_out           => s_data_out(43,45),
			out1               => s_out1(43,45),
			out2               => s_out2(43,45),
			lock_lower_row_out => s_locks_lower_out(43,45),
			lock_lower_row_in  => s_locks_lower_in(43,45),
			in1                => s_in1(43,45),
			in2                => s_in2(43,45),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(45)
		);
	s_in1(43,45)            <= s_out1(44,45);
	s_in2(43,45)            <= s_out2(44,46);
	s_locks_lower_in(43,45) <= s_locks_lower_out(44,45);

		normal_cell_43_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,46),
			fetch              => s_fetch(43,46),
			data_in            => s_data_in(43,46),
			data_out           => s_data_out(43,46),
			out1               => s_out1(43,46),
			out2               => s_out2(43,46),
			lock_lower_row_out => s_locks_lower_out(43,46),
			lock_lower_row_in  => s_locks_lower_in(43,46),
			in1                => s_in1(43,46),
			in2                => s_in2(43,46),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(46)
		);
	s_in1(43,46)            <= s_out1(44,46);
	s_in2(43,46)            <= s_out2(44,47);
	s_locks_lower_in(43,46) <= s_locks_lower_out(44,46);

		normal_cell_43_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,47),
			fetch              => s_fetch(43,47),
			data_in            => s_data_in(43,47),
			data_out           => s_data_out(43,47),
			out1               => s_out1(43,47),
			out2               => s_out2(43,47),
			lock_lower_row_out => s_locks_lower_out(43,47),
			lock_lower_row_in  => s_locks_lower_in(43,47),
			in1                => s_in1(43,47),
			in2                => s_in2(43,47),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(47)
		);
	s_in1(43,47)            <= s_out1(44,47);
	s_in2(43,47)            <= s_out2(44,48);
	s_locks_lower_in(43,47) <= s_locks_lower_out(44,47);

		normal_cell_43_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,48),
			fetch              => s_fetch(43,48),
			data_in            => s_data_in(43,48),
			data_out           => s_data_out(43,48),
			out1               => s_out1(43,48),
			out2               => s_out2(43,48),
			lock_lower_row_out => s_locks_lower_out(43,48),
			lock_lower_row_in  => s_locks_lower_in(43,48),
			in1                => s_in1(43,48),
			in2                => s_in2(43,48),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(48)
		);
	s_in1(43,48)            <= s_out1(44,48);
	s_in2(43,48)            <= s_out2(44,49);
	s_locks_lower_in(43,48) <= s_locks_lower_out(44,48);

		normal_cell_43_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,49),
			fetch              => s_fetch(43,49),
			data_in            => s_data_in(43,49),
			data_out           => s_data_out(43,49),
			out1               => s_out1(43,49),
			out2               => s_out2(43,49),
			lock_lower_row_out => s_locks_lower_out(43,49),
			lock_lower_row_in  => s_locks_lower_in(43,49),
			in1                => s_in1(43,49),
			in2                => s_in2(43,49),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(49)
		);
	s_in1(43,49)            <= s_out1(44,49);
	s_in2(43,49)            <= s_out2(44,50);
	s_locks_lower_in(43,49) <= s_locks_lower_out(44,49);

		normal_cell_43_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,50),
			fetch              => s_fetch(43,50),
			data_in            => s_data_in(43,50),
			data_out           => s_data_out(43,50),
			out1               => s_out1(43,50),
			out2               => s_out2(43,50),
			lock_lower_row_out => s_locks_lower_out(43,50),
			lock_lower_row_in  => s_locks_lower_in(43,50),
			in1                => s_in1(43,50),
			in2                => s_in2(43,50),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(50)
		);
	s_in1(43,50)            <= s_out1(44,50);
	s_in2(43,50)            <= s_out2(44,51);
	s_locks_lower_in(43,50) <= s_locks_lower_out(44,50);

		normal_cell_43_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,51),
			fetch              => s_fetch(43,51),
			data_in            => s_data_in(43,51),
			data_out           => s_data_out(43,51),
			out1               => s_out1(43,51),
			out2               => s_out2(43,51),
			lock_lower_row_out => s_locks_lower_out(43,51),
			lock_lower_row_in  => s_locks_lower_in(43,51),
			in1                => s_in1(43,51),
			in2                => s_in2(43,51),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(51)
		);
	s_in1(43,51)            <= s_out1(44,51);
	s_in2(43,51)            <= s_out2(44,52);
	s_locks_lower_in(43,51) <= s_locks_lower_out(44,51);

		normal_cell_43_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,52),
			fetch              => s_fetch(43,52),
			data_in            => s_data_in(43,52),
			data_out           => s_data_out(43,52),
			out1               => s_out1(43,52),
			out2               => s_out2(43,52),
			lock_lower_row_out => s_locks_lower_out(43,52),
			lock_lower_row_in  => s_locks_lower_in(43,52),
			in1                => s_in1(43,52),
			in2                => s_in2(43,52),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(52)
		);
	s_in1(43,52)            <= s_out1(44,52);
	s_in2(43,52)            <= s_out2(44,53);
	s_locks_lower_in(43,52) <= s_locks_lower_out(44,52);

		normal_cell_43_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,53),
			fetch              => s_fetch(43,53),
			data_in            => s_data_in(43,53),
			data_out           => s_data_out(43,53),
			out1               => s_out1(43,53),
			out2               => s_out2(43,53),
			lock_lower_row_out => s_locks_lower_out(43,53),
			lock_lower_row_in  => s_locks_lower_in(43,53),
			in1                => s_in1(43,53),
			in2                => s_in2(43,53),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(53)
		);
	s_in1(43,53)            <= s_out1(44,53);
	s_in2(43,53)            <= s_out2(44,54);
	s_locks_lower_in(43,53) <= s_locks_lower_out(44,53);

		normal_cell_43_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,54),
			fetch              => s_fetch(43,54),
			data_in            => s_data_in(43,54),
			data_out           => s_data_out(43,54),
			out1               => s_out1(43,54),
			out2               => s_out2(43,54),
			lock_lower_row_out => s_locks_lower_out(43,54),
			lock_lower_row_in  => s_locks_lower_in(43,54),
			in1                => s_in1(43,54),
			in2                => s_in2(43,54),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(54)
		);
	s_in1(43,54)            <= s_out1(44,54);
	s_in2(43,54)            <= s_out2(44,55);
	s_locks_lower_in(43,54) <= s_locks_lower_out(44,54);

		normal_cell_43_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,55),
			fetch              => s_fetch(43,55),
			data_in            => s_data_in(43,55),
			data_out           => s_data_out(43,55),
			out1               => s_out1(43,55),
			out2               => s_out2(43,55),
			lock_lower_row_out => s_locks_lower_out(43,55),
			lock_lower_row_in  => s_locks_lower_in(43,55),
			in1                => s_in1(43,55),
			in2                => s_in2(43,55),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(55)
		);
	s_in1(43,55)            <= s_out1(44,55);
	s_in2(43,55)            <= s_out2(44,56);
	s_locks_lower_in(43,55) <= s_locks_lower_out(44,55);

		normal_cell_43_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,56),
			fetch              => s_fetch(43,56),
			data_in            => s_data_in(43,56),
			data_out           => s_data_out(43,56),
			out1               => s_out1(43,56),
			out2               => s_out2(43,56),
			lock_lower_row_out => s_locks_lower_out(43,56),
			lock_lower_row_in  => s_locks_lower_in(43,56),
			in1                => s_in1(43,56),
			in2                => s_in2(43,56),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(56)
		);
	s_in1(43,56)            <= s_out1(44,56);
	s_in2(43,56)            <= s_out2(44,57);
	s_locks_lower_in(43,56) <= s_locks_lower_out(44,56);

		normal_cell_43_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,57),
			fetch              => s_fetch(43,57),
			data_in            => s_data_in(43,57),
			data_out           => s_data_out(43,57),
			out1               => s_out1(43,57),
			out2               => s_out2(43,57),
			lock_lower_row_out => s_locks_lower_out(43,57),
			lock_lower_row_in  => s_locks_lower_in(43,57),
			in1                => s_in1(43,57),
			in2                => s_in2(43,57),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(57)
		);
	s_in1(43,57)            <= s_out1(44,57);
	s_in2(43,57)            <= s_out2(44,58);
	s_locks_lower_in(43,57) <= s_locks_lower_out(44,57);

		normal_cell_43_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,58),
			fetch              => s_fetch(43,58),
			data_in            => s_data_in(43,58),
			data_out           => s_data_out(43,58),
			out1               => s_out1(43,58),
			out2               => s_out2(43,58),
			lock_lower_row_out => s_locks_lower_out(43,58),
			lock_lower_row_in  => s_locks_lower_in(43,58),
			in1                => s_in1(43,58),
			in2                => s_in2(43,58),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(58)
		);
	s_in1(43,58)            <= s_out1(44,58);
	s_in2(43,58)            <= s_out2(44,59);
	s_locks_lower_in(43,58) <= s_locks_lower_out(44,58);

		normal_cell_43_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,59),
			fetch              => s_fetch(43,59),
			data_in            => s_data_in(43,59),
			data_out           => s_data_out(43,59),
			out1               => s_out1(43,59),
			out2               => s_out2(43,59),
			lock_lower_row_out => s_locks_lower_out(43,59),
			lock_lower_row_in  => s_locks_lower_in(43,59),
			in1                => s_in1(43,59),
			in2                => s_in2(43,59),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(59)
		);
	s_in1(43,59)            <= s_out1(44,59);
	s_in2(43,59)            <= s_out2(44,60);
	s_locks_lower_in(43,59) <= s_locks_lower_out(44,59);

		last_col_cell_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(43,60),
			fetch              => s_fetch(43,60),
			data_in            => s_data_in(43,60),
			data_out           => s_data_out(43,60),
			out1               => s_out1(43,60),
			out2               => s_out2(43,60),
			lock_lower_row_out => s_locks_lower_out(43,60),
			lock_lower_row_in  => s_locks_lower_in(43,60),
			in1                => s_in1(43,60),
			in2                => (others => '0'),
			lock_row           => s_locks(43),
			piv_found          => s_piv_found,
			row_data           => s_row_data(43),
			col_data           => s_col_data(60)
		);
	s_in1(43,60)            <= s_out1(44,60);
	s_locks_lower_in(43,60) <= s_locks_lower_out(44,60);

		normal_cell_44_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,1),
			fetch              => s_fetch(44,1),
			data_in            => s_data_in(44,1),
			data_out           => s_data_out(44,1),
			out1               => s_out1(44,1),
			out2               => s_out2(44,1),
			lock_lower_row_out => s_locks_lower_out(44,1),
			lock_lower_row_in  => s_locks_lower_in(44,1),
			in1                => s_in1(44,1),
			in2                => s_in2(44,1),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(1)
		);
	s_in1(44,1)            <= s_out1(45,1);
	s_in2(44,1)            <= s_out2(45,2);
	s_locks_lower_in(44,1) <= s_locks_lower_out(45,1);

		normal_cell_44_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,2),
			fetch              => s_fetch(44,2),
			data_in            => s_data_in(44,2),
			data_out           => s_data_out(44,2),
			out1               => s_out1(44,2),
			out2               => s_out2(44,2),
			lock_lower_row_out => s_locks_lower_out(44,2),
			lock_lower_row_in  => s_locks_lower_in(44,2),
			in1                => s_in1(44,2),
			in2                => s_in2(44,2),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(2)
		);
	s_in1(44,2)            <= s_out1(45,2);
	s_in2(44,2)            <= s_out2(45,3);
	s_locks_lower_in(44,2) <= s_locks_lower_out(45,2);

		normal_cell_44_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,3),
			fetch              => s_fetch(44,3),
			data_in            => s_data_in(44,3),
			data_out           => s_data_out(44,3),
			out1               => s_out1(44,3),
			out2               => s_out2(44,3),
			lock_lower_row_out => s_locks_lower_out(44,3),
			lock_lower_row_in  => s_locks_lower_in(44,3),
			in1                => s_in1(44,3),
			in2                => s_in2(44,3),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(3)
		);
	s_in1(44,3)            <= s_out1(45,3);
	s_in2(44,3)            <= s_out2(45,4);
	s_locks_lower_in(44,3) <= s_locks_lower_out(45,3);

		normal_cell_44_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,4),
			fetch              => s_fetch(44,4),
			data_in            => s_data_in(44,4),
			data_out           => s_data_out(44,4),
			out1               => s_out1(44,4),
			out2               => s_out2(44,4),
			lock_lower_row_out => s_locks_lower_out(44,4),
			lock_lower_row_in  => s_locks_lower_in(44,4),
			in1                => s_in1(44,4),
			in2                => s_in2(44,4),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(4)
		);
	s_in1(44,4)            <= s_out1(45,4);
	s_in2(44,4)            <= s_out2(45,5);
	s_locks_lower_in(44,4) <= s_locks_lower_out(45,4);

		normal_cell_44_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,5),
			fetch              => s_fetch(44,5),
			data_in            => s_data_in(44,5),
			data_out           => s_data_out(44,5),
			out1               => s_out1(44,5),
			out2               => s_out2(44,5),
			lock_lower_row_out => s_locks_lower_out(44,5),
			lock_lower_row_in  => s_locks_lower_in(44,5),
			in1                => s_in1(44,5),
			in2                => s_in2(44,5),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(5)
		);
	s_in1(44,5)            <= s_out1(45,5);
	s_in2(44,5)            <= s_out2(45,6);
	s_locks_lower_in(44,5) <= s_locks_lower_out(45,5);

		normal_cell_44_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,6),
			fetch              => s_fetch(44,6),
			data_in            => s_data_in(44,6),
			data_out           => s_data_out(44,6),
			out1               => s_out1(44,6),
			out2               => s_out2(44,6),
			lock_lower_row_out => s_locks_lower_out(44,6),
			lock_lower_row_in  => s_locks_lower_in(44,6),
			in1                => s_in1(44,6),
			in2                => s_in2(44,6),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(6)
		);
	s_in1(44,6)            <= s_out1(45,6);
	s_in2(44,6)            <= s_out2(45,7);
	s_locks_lower_in(44,6) <= s_locks_lower_out(45,6);

		normal_cell_44_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,7),
			fetch              => s_fetch(44,7),
			data_in            => s_data_in(44,7),
			data_out           => s_data_out(44,7),
			out1               => s_out1(44,7),
			out2               => s_out2(44,7),
			lock_lower_row_out => s_locks_lower_out(44,7),
			lock_lower_row_in  => s_locks_lower_in(44,7),
			in1                => s_in1(44,7),
			in2                => s_in2(44,7),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(7)
		);
	s_in1(44,7)            <= s_out1(45,7);
	s_in2(44,7)            <= s_out2(45,8);
	s_locks_lower_in(44,7) <= s_locks_lower_out(45,7);

		normal_cell_44_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,8),
			fetch              => s_fetch(44,8),
			data_in            => s_data_in(44,8),
			data_out           => s_data_out(44,8),
			out1               => s_out1(44,8),
			out2               => s_out2(44,8),
			lock_lower_row_out => s_locks_lower_out(44,8),
			lock_lower_row_in  => s_locks_lower_in(44,8),
			in1                => s_in1(44,8),
			in2                => s_in2(44,8),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(8)
		);
	s_in1(44,8)            <= s_out1(45,8);
	s_in2(44,8)            <= s_out2(45,9);
	s_locks_lower_in(44,8) <= s_locks_lower_out(45,8);

		normal_cell_44_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,9),
			fetch              => s_fetch(44,9),
			data_in            => s_data_in(44,9),
			data_out           => s_data_out(44,9),
			out1               => s_out1(44,9),
			out2               => s_out2(44,9),
			lock_lower_row_out => s_locks_lower_out(44,9),
			lock_lower_row_in  => s_locks_lower_in(44,9),
			in1                => s_in1(44,9),
			in2                => s_in2(44,9),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(9)
		);
	s_in1(44,9)            <= s_out1(45,9);
	s_in2(44,9)            <= s_out2(45,10);
	s_locks_lower_in(44,9) <= s_locks_lower_out(45,9);

		normal_cell_44_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,10),
			fetch              => s_fetch(44,10),
			data_in            => s_data_in(44,10),
			data_out           => s_data_out(44,10),
			out1               => s_out1(44,10),
			out2               => s_out2(44,10),
			lock_lower_row_out => s_locks_lower_out(44,10),
			lock_lower_row_in  => s_locks_lower_in(44,10),
			in1                => s_in1(44,10),
			in2                => s_in2(44,10),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(10)
		);
	s_in1(44,10)            <= s_out1(45,10);
	s_in2(44,10)            <= s_out2(45,11);
	s_locks_lower_in(44,10) <= s_locks_lower_out(45,10);

		normal_cell_44_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,11),
			fetch              => s_fetch(44,11),
			data_in            => s_data_in(44,11),
			data_out           => s_data_out(44,11),
			out1               => s_out1(44,11),
			out2               => s_out2(44,11),
			lock_lower_row_out => s_locks_lower_out(44,11),
			lock_lower_row_in  => s_locks_lower_in(44,11),
			in1                => s_in1(44,11),
			in2                => s_in2(44,11),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(11)
		);
	s_in1(44,11)            <= s_out1(45,11);
	s_in2(44,11)            <= s_out2(45,12);
	s_locks_lower_in(44,11) <= s_locks_lower_out(45,11);

		normal_cell_44_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,12),
			fetch              => s_fetch(44,12),
			data_in            => s_data_in(44,12),
			data_out           => s_data_out(44,12),
			out1               => s_out1(44,12),
			out2               => s_out2(44,12),
			lock_lower_row_out => s_locks_lower_out(44,12),
			lock_lower_row_in  => s_locks_lower_in(44,12),
			in1                => s_in1(44,12),
			in2                => s_in2(44,12),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(12)
		);
	s_in1(44,12)            <= s_out1(45,12);
	s_in2(44,12)            <= s_out2(45,13);
	s_locks_lower_in(44,12) <= s_locks_lower_out(45,12);

		normal_cell_44_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,13),
			fetch              => s_fetch(44,13),
			data_in            => s_data_in(44,13),
			data_out           => s_data_out(44,13),
			out1               => s_out1(44,13),
			out2               => s_out2(44,13),
			lock_lower_row_out => s_locks_lower_out(44,13),
			lock_lower_row_in  => s_locks_lower_in(44,13),
			in1                => s_in1(44,13),
			in2                => s_in2(44,13),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(13)
		);
	s_in1(44,13)            <= s_out1(45,13);
	s_in2(44,13)            <= s_out2(45,14);
	s_locks_lower_in(44,13) <= s_locks_lower_out(45,13);

		normal_cell_44_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,14),
			fetch              => s_fetch(44,14),
			data_in            => s_data_in(44,14),
			data_out           => s_data_out(44,14),
			out1               => s_out1(44,14),
			out2               => s_out2(44,14),
			lock_lower_row_out => s_locks_lower_out(44,14),
			lock_lower_row_in  => s_locks_lower_in(44,14),
			in1                => s_in1(44,14),
			in2                => s_in2(44,14),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(14)
		);
	s_in1(44,14)            <= s_out1(45,14);
	s_in2(44,14)            <= s_out2(45,15);
	s_locks_lower_in(44,14) <= s_locks_lower_out(45,14);

		normal_cell_44_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,15),
			fetch              => s_fetch(44,15),
			data_in            => s_data_in(44,15),
			data_out           => s_data_out(44,15),
			out1               => s_out1(44,15),
			out2               => s_out2(44,15),
			lock_lower_row_out => s_locks_lower_out(44,15),
			lock_lower_row_in  => s_locks_lower_in(44,15),
			in1                => s_in1(44,15),
			in2                => s_in2(44,15),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(15)
		);
	s_in1(44,15)            <= s_out1(45,15);
	s_in2(44,15)            <= s_out2(45,16);
	s_locks_lower_in(44,15) <= s_locks_lower_out(45,15);

		normal_cell_44_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,16),
			fetch              => s_fetch(44,16),
			data_in            => s_data_in(44,16),
			data_out           => s_data_out(44,16),
			out1               => s_out1(44,16),
			out2               => s_out2(44,16),
			lock_lower_row_out => s_locks_lower_out(44,16),
			lock_lower_row_in  => s_locks_lower_in(44,16),
			in1                => s_in1(44,16),
			in2                => s_in2(44,16),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(16)
		);
	s_in1(44,16)            <= s_out1(45,16);
	s_in2(44,16)            <= s_out2(45,17);
	s_locks_lower_in(44,16) <= s_locks_lower_out(45,16);

		normal_cell_44_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,17),
			fetch              => s_fetch(44,17),
			data_in            => s_data_in(44,17),
			data_out           => s_data_out(44,17),
			out1               => s_out1(44,17),
			out2               => s_out2(44,17),
			lock_lower_row_out => s_locks_lower_out(44,17),
			lock_lower_row_in  => s_locks_lower_in(44,17),
			in1                => s_in1(44,17),
			in2                => s_in2(44,17),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(17)
		);
	s_in1(44,17)            <= s_out1(45,17);
	s_in2(44,17)            <= s_out2(45,18);
	s_locks_lower_in(44,17) <= s_locks_lower_out(45,17);

		normal_cell_44_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,18),
			fetch              => s_fetch(44,18),
			data_in            => s_data_in(44,18),
			data_out           => s_data_out(44,18),
			out1               => s_out1(44,18),
			out2               => s_out2(44,18),
			lock_lower_row_out => s_locks_lower_out(44,18),
			lock_lower_row_in  => s_locks_lower_in(44,18),
			in1                => s_in1(44,18),
			in2                => s_in2(44,18),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(18)
		);
	s_in1(44,18)            <= s_out1(45,18);
	s_in2(44,18)            <= s_out2(45,19);
	s_locks_lower_in(44,18) <= s_locks_lower_out(45,18);

		normal_cell_44_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,19),
			fetch              => s_fetch(44,19),
			data_in            => s_data_in(44,19),
			data_out           => s_data_out(44,19),
			out1               => s_out1(44,19),
			out2               => s_out2(44,19),
			lock_lower_row_out => s_locks_lower_out(44,19),
			lock_lower_row_in  => s_locks_lower_in(44,19),
			in1                => s_in1(44,19),
			in2                => s_in2(44,19),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(19)
		);
	s_in1(44,19)            <= s_out1(45,19);
	s_in2(44,19)            <= s_out2(45,20);
	s_locks_lower_in(44,19) <= s_locks_lower_out(45,19);

		normal_cell_44_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,20),
			fetch              => s_fetch(44,20),
			data_in            => s_data_in(44,20),
			data_out           => s_data_out(44,20),
			out1               => s_out1(44,20),
			out2               => s_out2(44,20),
			lock_lower_row_out => s_locks_lower_out(44,20),
			lock_lower_row_in  => s_locks_lower_in(44,20),
			in1                => s_in1(44,20),
			in2                => s_in2(44,20),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(20)
		);
	s_in1(44,20)            <= s_out1(45,20);
	s_in2(44,20)            <= s_out2(45,21);
	s_locks_lower_in(44,20) <= s_locks_lower_out(45,20);

		normal_cell_44_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,21),
			fetch              => s_fetch(44,21),
			data_in            => s_data_in(44,21),
			data_out           => s_data_out(44,21),
			out1               => s_out1(44,21),
			out2               => s_out2(44,21),
			lock_lower_row_out => s_locks_lower_out(44,21),
			lock_lower_row_in  => s_locks_lower_in(44,21),
			in1                => s_in1(44,21),
			in2                => s_in2(44,21),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(21)
		);
	s_in1(44,21)            <= s_out1(45,21);
	s_in2(44,21)            <= s_out2(45,22);
	s_locks_lower_in(44,21) <= s_locks_lower_out(45,21);

		normal_cell_44_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,22),
			fetch              => s_fetch(44,22),
			data_in            => s_data_in(44,22),
			data_out           => s_data_out(44,22),
			out1               => s_out1(44,22),
			out2               => s_out2(44,22),
			lock_lower_row_out => s_locks_lower_out(44,22),
			lock_lower_row_in  => s_locks_lower_in(44,22),
			in1                => s_in1(44,22),
			in2                => s_in2(44,22),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(22)
		);
	s_in1(44,22)            <= s_out1(45,22);
	s_in2(44,22)            <= s_out2(45,23);
	s_locks_lower_in(44,22) <= s_locks_lower_out(45,22);

		normal_cell_44_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,23),
			fetch              => s_fetch(44,23),
			data_in            => s_data_in(44,23),
			data_out           => s_data_out(44,23),
			out1               => s_out1(44,23),
			out2               => s_out2(44,23),
			lock_lower_row_out => s_locks_lower_out(44,23),
			lock_lower_row_in  => s_locks_lower_in(44,23),
			in1                => s_in1(44,23),
			in2                => s_in2(44,23),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(23)
		);
	s_in1(44,23)            <= s_out1(45,23);
	s_in2(44,23)            <= s_out2(45,24);
	s_locks_lower_in(44,23) <= s_locks_lower_out(45,23);

		normal_cell_44_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,24),
			fetch              => s_fetch(44,24),
			data_in            => s_data_in(44,24),
			data_out           => s_data_out(44,24),
			out1               => s_out1(44,24),
			out2               => s_out2(44,24),
			lock_lower_row_out => s_locks_lower_out(44,24),
			lock_lower_row_in  => s_locks_lower_in(44,24),
			in1                => s_in1(44,24),
			in2                => s_in2(44,24),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(24)
		);
	s_in1(44,24)            <= s_out1(45,24);
	s_in2(44,24)            <= s_out2(45,25);
	s_locks_lower_in(44,24) <= s_locks_lower_out(45,24);

		normal_cell_44_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,25),
			fetch              => s_fetch(44,25),
			data_in            => s_data_in(44,25),
			data_out           => s_data_out(44,25),
			out1               => s_out1(44,25),
			out2               => s_out2(44,25),
			lock_lower_row_out => s_locks_lower_out(44,25),
			lock_lower_row_in  => s_locks_lower_in(44,25),
			in1                => s_in1(44,25),
			in2                => s_in2(44,25),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(25)
		);
	s_in1(44,25)            <= s_out1(45,25);
	s_in2(44,25)            <= s_out2(45,26);
	s_locks_lower_in(44,25) <= s_locks_lower_out(45,25);

		normal_cell_44_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,26),
			fetch              => s_fetch(44,26),
			data_in            => s_data_in(44,26),
			data_out           => s_data_out(44,26),
			out1               => s_out1(44,26),
			out2               => s_out2(44,26),
			lock_lower_row_out => s_locks_lower_out(44,26),
			lock_lower_row_in  => s_locks_lower_in(44,26),
			in1                => s_in1(44,26),
			in2                => s_in2(44,26),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(26)
		);
	s_in1(44,26)            <= s_out1(45,26);
	s_in2(44,26)            <= s_out2(45,27);
	s_locks_lower_in(44,26) <= s_locks_lower_out(45,26);

		normal_cell_44_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,27),
			fetch              => s_fetch(44,27),
			data_in            => s_data_in(44,27),
			data_out           => s_data_out(44,27),
			out1               => s_out1(44,27),
			out2               => s_out2(44,27),
			lock_lower_row_out => s_locks_lower_out(44,27),
			lock_lower_row_in  => s_locks_lower_in(44,27),
			in1                => s_in1(44,27),
			in2                => s_in2(44,27),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(27)
		);
	s_in1(44,27)            <= s_out1(45,27);
	s_in2(44,27)            <= s_out2(45,28);
	s_locks_lower_in(44,27) <= s_locks_lower_out(45,27);

		normal_cell_44_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,28),
			fetch              => s_fetch(44,28),
			data_in            => s_data_in(44,28),
			data_out           => s_data_out(44,28),
			out1               => s_out1(44,28),
			out2               => s_out2(44,28),
			lock_lower_row_out => s_locks_lower_out(44,28),
			lock_lower_row_in  => s_locks_lower_in(44,28),
			in1                => s_in1(44,28),
			in2                => s_in2(44,28),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(28)
		);
	s_in1(44,28)            <= s_out1(45,28);
	s_in2(44,28)            <= s_out2(45,29);
	s_locks_lower_in(44,28) <= s_locks_lower_out(45,28);

		normal_cell_44_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,29),
			fetch              => s_fetch(44,29),
			data_in            => s_data_in(44,29),
			data_out           => s_data_out(44,29),
			out1               => s_out1(44,29),
			out2               => s_out2(44,29),
			lock_lower_row_out => s_locks_lower_out(44,29),
			lock_lower_row_in  => s_locks_lower_in(44,29),
			in1                => s_in1(44,29),
			in2                => s_in2(44,29),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(29)
		);
	s_in1(44,29)            <= s_out1(45,29);
	s_in2(44,29)            <= s_out2(45,30);
	s_locks_lower_in(44,29) <= s_locks_lower_out(45,29);

		normal_cell_44_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,30),
			fetch              => s_fetch(44,30),
			data_in            => s_data_in(44,30),
			data_out           => s_data_out(44,30),
			out1               => s_out1(44,30),
			out2               => s_out2(44,30),
			lock_lower_row_out => s_locks_lower_out(44,30),
			lock_lower_row_in  => s_locks_lower_in(44,30),
			in1                => s_in1(44,30),
			in2                => s_in2(44,30),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(30)
		);
	s_in1(44,30)            <= s_out1(45,30);
	s_in2(44,30)            <= s_out2(45,31);
	s_locks_lower_in(44,30) <= s_locks_lower_out(45,30);

		normal_cell_44_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,31),
			fetch              => s_fetch(44,31),
			data_in            => s_data_in(44,31),
			data_out           => s_data_out(44,31),
			out1               => s_out1(44,31),
			out2               => s_out2(44,31),
			lock_lower_row_out => s_locks_lower_out(44,31),
			lock_lower_row_in  => s_locks_lower_in(44,31),
			in1                => s_in1(44,31),
			in2                => s_in2(44,31),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(31)
		);
	s_in1(44,31)            <= s_out1(45,31);
	s_in2(44,31)            <= s_out2(45,32);
	s_locks_lower_in(44,31) <= s_locks_lower_out(45,31);

		normal_cell_44_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,32),
			fetch              => s_fetch(44,32),
			data_in            => s_data_in(44,32),
			data_out           => s_data_out(44,32),
			out1               => s_out1(44,32),
			out2               => s_out2(44,32),
			lock_lower_row_out => s_locks_lower_out(44,32),
			lock_lower_row_in  => s_locks_lower_in(44,32),
			in1                => s_in1(44,32),
			in2                => s_in2(44,32),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(32)
		);
	s_in1(44,32)            <= s_out1(45,32);
	s_in2(44,32)            <= s_out2(45,33);
	s_locks_lower_in(44,32) <= s_locks_lower_out(45,32);

		normal_cell_44_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,33),
			fetch              => s_fetch(44,33),
			data_in            => s_data_in(44,33),
			data_out           => s_data_out(44,33),
			out1               => s_out1(44,33),
			out2               => s_out2(44,33),
			lock_lower_row_out => s_locks_lower_out(44,33),
			lock_lower_row_in  => s_locks_lower_in(44,33),
			in1                => s_in1(44,33),
			in2                => s_in2(44,33),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(33)
		);
	s_in1(44,33)            <= s_out1(45,33);
	s_in2(44,33)            <= s_out2(45,34);
	s_locks_lower_in(44,33) <= s_locks_lower_out(45,33);

		normal_cell_44_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,34),
			fetch              => s_fetch(44,34),
			data_in            => s_data_in(44,34),
			data_out           => s_data_out(44,34),
			out1               => s_out1(44,34),
			out2               => s_out2(44,34),
			lock_lower_row_out => s_locks_lower_out(44,34),
			lock_lower_row_in  => s_locks_lower_in(44,34),
			in1                => s_in1(44,34),
			in2                => s_in2(44,34),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(34)
		);
	s_in1(44,34)            <= s_out1(45,34);
	s_in2(44,34)            <= s_out2(45,35);
	s_locks_lower_in(44,34) <= s_locks_lower_out(45,34);

		normal_cell_44_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,35),
			fetch              => s_fetch(44,35),
			data_in            => s_data_in(44,35),
			data_out           => s_data_out(44,35),
			out1               => s_out1(44,35),
			out2               => s_out2(44,35),
			lock_lower_row_out => s_locks_lower_out(44,35),
			lock_lower_row_in  => s_locks_lower_in(44,35),
			in1                => s_in1(44,35),
			in2                => s_in2(44,35),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(35)
		);
	s_in1(44,35)            <= s_out1(45,35);
	s_in2(44,35)            <= s_out2(45,36);
	s_locks_lower_in(44,35) <= s_locks_lower_out(45,35);

		normal_cell_44_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,36),
			fetch              => s_fetch(44,36),
			data_in            => s_data_in(44,36),
			data_out           => s_data_out(44,36),
			out1               => s_out1(44,36),
			out2               => s_out2(44,36),
			lock_lower_row_out => s_locks_lower_out(44,36),
			lock_lower_row_in  => s_locks_lower_in(44,36),
			in1                => s_in1(44,36),
			in2                => s_in2(44,36),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(36)
		);
	s_in1(44,36)            <= s_out1(45,36);
	s_in2(44,36)            <= s_out2(45,37);
	s_locks_lower_in(44,36) <= s_locks_lower_out(45,36);

		normal_cell_44_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,37),
			fetch              => s_fetch(44,37),
			data_in            => s_data_in(44,37),
			data_out           => s_data_out(44,37),
			out1               => s_out1(44,37),
			out2               => s_out2(44,37),
			lock_lower_row_out => s_locks_lower_out(44,37),
			lock_lower_row_in  => s_locks_lower_in(44,37),
			in1                => s_in1(44,37),
			in2                => s_in2(44,37),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(37)
		);
	s_in1(44,37)            <= s_out1(45,37);
	s_in2(44,37)            <= s_out2(45,38);
	s_locks_lower_in(44,37) <= s_locks_lower_out(45,37);

		normal_cell_44_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,38),
			fetch              => s_fetch(44,38),
			data_in            => s_data_in(44,38),
			data_out           => s_data_out(44,38),
			out1               => s_out1(44,38),
			out2               => s_out2(44,38),
			lock_lower_row_out => s_locks_lower_out(44,38),
			lock_lower_row_in  => s_locks_lower_in(44,38),
			in1                => s_in1(44,38),
			in2                => s_in2(44,38),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(38)
		);
	s_in1(44,38)            <= s_out1(45,38);
	s_in2(44,38)            <= s_out2(45,39);
	s_locks_lower_in(44,38) <= s_locks_lower_out(45,38);

		normal_cell_44_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,39),
			fetch              => s_fetch(44,39),
			data_in            => s_data_in(44,39),
			data_out           => s_data_out(44,39),
			out1               => s_out1(44,39),
			out2               => s_out2(44,39),
			lock_lower_row_out => s_locks_lower_out(44,39),
			lock_lower_row_in  => s_locks_lower_in(44,39),
			in1                => s_in1(44,39),
			in2                => s_in2(44,39),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(39)
		);
	s_in1(44,39)            <= s_out1(45,39);
	s_in2(44,39)            <= s_out2(45,40);
	s_locks_lower_in(44,39) <= s_locks_lower_out(45,39);

		normal_cell_44_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,40),
			fetch              => s_fetch(44,40),
			data_in            => s_data_in(44,40),
			data_out           => s_data_out(44,40),
			out1               => s_out1(44,40),
			out2               => s_out2(44,40),
			lock_lower_row_out => s_locks_lower_out(44,40),
			lock_lower_row_in  => s_locks_lower_in(44,40),
			in1                => s_in1(44,40),
			in2                => s_in2(44,40),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(40)
		);
	s_in1(44,40)            <= s_out1(45,40);
	s_in2(44,40)            <= s_out2(45,41);
	s_locks_lower_in(44,40) <= s_locks_lower_out(45,40);

		normal_cell_44_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,41),
			fetch              => s_fetch(44,41),
			data_in            => s_data_in(44,41),
			data_out           => s_data_out(44,41),
			out1               => s_out1(44,41),
			out2               => s_out2(44,41),
			lock_lower_row_out => s_locks_lower_out(44,41),
			lock_lower_row_in  => s_locks_lower_in(44,41),
			in1                => s_in1(44,41),
			in2                => s_in2(44,41),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(41)
		);
	s_in1(44,41)            <= s_out1(45,41);
	s_in2(44,41)            <= s_out2(45,42);
	s_locks_lower_in(44,41) <= s_locks_lower_out(45,41);

		normal_cell_44_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,42),
			fetch              => s_fetch(44,42),
			data_in            => s_data_in(44,42),
			data_out           => s_data_out(44,42),
			out1               => s_out1(44,42),
			out2               => s_out2(44,42),
			lock_lower_row_out => s_locks_lower_out(44,42),
			lock_lower_row_in  => s_locks_lower_in(44,42),
			in1                => s_in1(44,42),
			in2                => s_in2(44,42),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(42)
		);
	s_in1(44,42)            <= s_out1(45,42);
	s_in2(44,42)            <= s_out2(45,43);
	s_locks_lower_in(44,42) <= s_locks_lower_out(45,42);

		normal_cell_44_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,43),
			fetch              => s_fetch(44,43),
			data_in            => s_data_in(44,43),
			data_out           => s_data_out(44,43),
			out1               => s_out1(44,43),
			out2               => s_out2(44,43),
			lock_lower_row_out => s_locks_lower_out(44,43),
			lock_lower_row_in  => s_locks_lower_in(44,43),
			in1                => s_in1(44,43),
			in2                => s_in2(44,43),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(43)
		);
	s_in1(44,43)            <= s_out1(45,43);
	s_in2(44,43)            <= s_out2(45,44);
	s_locks_lower_in(44,43) <= s_locks_lower_out(45,43);

		normal_cell_44_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,44),
			fetch              => s_fetch(44,44),
			data_in            => s_data_in(44,44),
			data_out           => s_data_out(44,44),
			out1               => s_out1(44,44),
			out2               => s_out2(44,44),
			lock_lower_row_out => s_locks_lower_out(44,44),
			lock_lower_row_in  => s_locks_lower_in(44,44),
			in1                => s_in1(44,44),
			in2                => s_in2(44,44),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(44)
		);
	s_in1(44,44)            <= s_out1(45,44);
	s_in2(44,44)            <= s_out2(45,45);
	s_locks_lower_in(44,44) <= s_locks_lower_out(45,44);

		normal_cell_44_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,45),
			fetch              => s_fetch(44,45),
			data_in            => s_data_in(44,45),
			data_out           => s_data_out(44,45),
			out1               => s_out1(44,45),
			out2               => s_out2(44,45),
			lock_lower_row_out => s_locks_lower_out(44,45),
			lock_lower_row_in  => s_locks_lower_in(44,45),
			in1                => s_in1(44,45),
			in2                => s_in2(44,45),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(45)
		);
	s_in1(44,45)            <= s_out1(45,45);
	s_in2(44,45)            <= s_out2(45,46);
	s_locks_lower_in(44,45) <= s_locks_lower_out(45,45);

		normal_cell_44_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,46),
			fetch              => s_fetch(44,46),
			data_in            => s_data_in(44,46),
			data_out           => s_data_out(44,46),
			out1               => s_out1(44,46),
			out2               => s_out2(44,46),
			lock_lower_row_out => s_locks_lower_out(44,46),
			lock_lower_row_in  => s_locks_lower_in(44,46),
			in1                => s_in1(44,46),
			in2                => s_in2(44,46),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(46)
		);
	s_in1(44,46)            <= s_out1(45,46);
	s_in2(44,46)            <= s_out2(45,47);
	s_locks_lower_in(44,46) <= s_locks_lower_out(45,46);

		normal_cell_44_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,47),
			fetch              => s_fetch(44,47),
			data_in            => s_data_in(44,47),
			data_out           => s_data_out(44,47),
			out1               => s_out1(44,47),
			out2               => s_out2(44,47),
			lock_lower_row_out => s_locks_lower_out(44,47),
			lock_lower_row_in  => s_locks_lower_in(44,47),
			in1                => s_in1(44,47),
			in2                => s_in2(44,47),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(47)
		);
	s_in1(44,47)            <= s_out1(45,47);
	s_in2(44,47)            <= s_out2(45,48);
	s_locks_lower_in(44,47) <= s_locks_lower_out(45,47);

		normal_cell_44_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,48),
			fetch              => s_fetch(44,48),
			data_in            => s_data_in(44,48),
			data_out           => s_data_out(44,48),
			out1               => s_out1(44,48),
			out2               => s_out2(44,48),
			lock_lower_row_out => s_locks_lower_out(44,48),
			lock_lower_row_in  => s_locks_lower_in(44,48),
			in1                => s_in1(44,48),
			in2                => s_in2(44,48),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(48)
		);
	s_in1(44,48)            <= s_out1(45,48);
	s_in2(44,48)            <= s_out2(45,49);
	s_locks_lower_in(44,48) <= s_locks_lower_out(45,48);

		normal_cell_44_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,49),
			fetch              => s_fetch(44,49),
			data_in            => s_data_in(44,49),
			data_out           => s_data_out(44,49),
			out1               => s_out1(44,49),
			out2               => s_out2(44,49),
			lock_lower_row_out => s_locks_lower_out(44,49),
			lock_lower_row_in  => s_locks_lower_in(44,49),
			in1                => s_in1(44,49),
			in2                => s_in2(44,49),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(49)
		);
	s_in1(44,49)            <= s_out1(45,49);
	s_in2(44,49)            <= s_out2(45,50);
	s_locks_lower_in(44,49) <= s_locks_lower_out(45,49);

		normal_cell_44_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,50),
			fetch              => s_fetch(44,50),
			data_in            => s_data_in(44,50),
			data_out           => s_data_out(44,50),
			out1               => s_out1(44,50),
			out2               => s_out2(44,50),
			lock_lower_row_out => s_locks_lower_out(44,50),
			lock_lower_row_in  => s_locks_lower_in(44,50),
			in1                => s_in1(44,50),
			in2                => s_in2(44,50),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(50)
		);
	s_in1(44,50)            <= s_out1(45,50);
	s_in2(44,50)            <= s_out2(45,51);
	s_locks_lower_in(44,50) <= s_locks_lower_out(45,50);

		normal_cell_44_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,51),
			fetch              => s_fetch(44,51),
			data_in            => s_data_in(44,51),
			data_out           => s_data_out(44,51),
			out1               => s_out1(44,51),
			out2               => s_out2(44,51),
			lock_lower_row_out => s_locks_lower_out(44,51),
			lock_lower_row_in  => s_locks_lower_in(44,51),
			in1                => s_in1(44,51),
			in2                => s_in2(44,51),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(51)
		);
	s_in1(44,51)            <= s_out1(45,51);
	s_in2(44,51)            <= s_out2(45,52);
	s_locks_lower_in(44,51) <= s_locks_lower_out(45,51);

		normal_cell_44_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,52),
			fetch              => s_fetch(44,52),
			data_in            => s_data_in(44,52),
			data_out           => s_data_out(44,52),
			out1               => s_out1(44,52),
			out2               => s_out2(44,52),
			lock_lower_row_out => s_locks_lower_out(44,52),
			lock_lower_row_in  => s_locks_lower_in(44,52),
			in1                => s_in1(44,52),
			in2                => s_in2(44,52),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(52)
		);
	s_in1(44,52)            <= s_out1(45,52);
	s_in2(44,52)            <= s_out2(45,53);
	s_locks_lower_in(44,52) <= s_locks_lower_out(45,52);

		normal_cell_44_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,53),
			fetch              => s_fetch(44,53),
			data_in            => s_data_in(44,53),
			data_out           => s_data_out(44,53),
			out1               => s_out1(44,53),
			out2               => s_out2(44,53),
			lock_lower_row_out => s_locks_lower_out(44,53),
			lock_lower_row_in  => s_locks_lower_in(44,53),
			in1                => s_in1(44,53),
			in2                => s_in2(44,53),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(53)
		);
	s_in1(44,53)            <= s_out1(45,53);
	s_in2(44,53)            <= s_out2(45,54);
	s_locks_lower_in(44,53) <= s_locks_lower_out(45,53);

		normal_cell_44_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,54),
			fetch              => s_fetch(44,54),
			data_in            => s_data_in(44,54),
			data_out           => s_data_out(44,54),
			out1               => s_out1(44,54),
			out2               => s_out2(44,54),
			lock_lower_row_out => s_locks_lower_out(44,54),
			lock_lower_row_in  => s_locks_lower_in(44,54),
			in1                => s_in1(44,54),
			in2                => s_in2(44,54),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(54)
		);
	s_in1(44,54)            <= s_out1(45,54);
	s_in2(44,54)            <= s_out2(45,55);
	s_locks_lower_in(44,54) <= s_locks_lower_out(45,54);

		normal_cell_44_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,55),
			fetch              => s_fetch(44,55),
			data_in            => s_data_in(44,55),
			data_out           => s_data_out(44,55),
			out1               => s_out1(44,55),
			out2               => s_out2(44,55),
			lock_lower_row_out => s_locks_lower_out(44,55),
			lock_lower_row_in  => s_locks_lower_in(44,55),
			in1                => s_in1(44,55),
			in2                => s_in2(44,55),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(55)
		);
	s_in1(44,55)            <= s_out1(45,55);
	s_in2(44,55)            <= s_out2(45,56);
	s_locks_lower_in(44,55) <= s_locks_lower_out(45,55);

		normal_cell_44_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,56),
			fetch              => s_fetch(44,56),
			data_in            => s_data_in(44,56),
			data_out           => s_data_out(44,56),
			out1               => s_out1(44,56),
			out2               => s_out2(44,56),
			lock_lower_row_out => s_locks_lower_out(44,56),
			lock_lower_row_in  => s_locks_lower_in(44,56),
			in1                => s_in1(44,56),
			in2                => s_in2(44,56),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(56)
		);
	s_in1(44,56)            <= s_out1(45,56);
	s_in2(44,56)            <= s_out2(45,57);
	s_locks_lower_in(44,56) <= s_locks_lower_out(45,56);

		normal_cell_44_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,57),
			fetch              => s_fetch(44,57),
			data_in            => s_data_in(44,57),
			data_out           => s_data_out(44,57),
			out1               => s_out1(44,57),
			out2               => s_out2(44,57),
			lock_lower_row_out => s_locks_lower_out(44,57),
			lock_lower_row_in  => s_locks_lower_in(44,57),
			in1                => s_in1(44,57),
			in2                => s_in2(44,57),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(57)
		);
	s_in1(44,57)            <= s_out1(45,57);
	s_in2(44,57)            <= s_out2(45,58);
	s_locks_lower_in(44,57) <= s_locks_lower_out(45,57);

		normal_cell_44_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,58),
			fetch              => s_fetch(44,58),
			data_in            => s_data_in(44,58),
			data_out           => s_data_out(44,58),
			out1               => s_out1(44,58),
			out2               => s_out2(44,58),
			lock_lower_row_out => s_locks_lower_out(44,58),
			lock_lower_row_in  => s_locks_lower_in(44,58),
			in1                => s_in1(44,58),
			in2                => s_in2(44,58),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(58)
		);
	s_in1(44,58)            <= s_out1(45,58);
	s_in2(44,58)            <= s_out2(45,59);
	s_locks_lower_in(44,58) <= s_locks_lower_out(45,58);

		normal_cell_44_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,59),
			fetch              => s_fetch(44,59),
			data_in            => s_data_in(44,59),
			data_out           => s_data_out(44,59),
			out1               => s_out1(44,59),
			out2               => s_out2(44,59),
			lock_lower_row_out => s_locks_lower_out(44,59),
			lock_lower_row_in  => s_locks_lower_in(44,59),
			in1                => s_in1(44,59),
			in2                => s_in2(44,59),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(59)
		);
	s_in1(44,59)            <= s_out1(45,59);
	s_in2(44,59)            <= s_out2(45,60);
	s_locks_lower_in(44,59) <= s_locks_lower_out(45,59);

		last_col_cell_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(44,60),
			fetch              => s_fetch(44,60),
			data_in            => s_data_in(44,60),
			data_out           => s_data_out(44,60),
			out1               => s_out1(44,60),
			out2               => s_out2(44,60),
			lock_lower_row_out => s_locks_lower_out(44,60),
			lock_lower_row_in  => s_locks_lower_in(44,60),
			in1                => s_in1(44,60),
			in2                => (others => '0'),
			lock_row           => s_locks(44),
			piv_found          => s_piv_found,
			row_data           => s_row_data(44),
			col_data           => s_col_data(60)
		);
	s_in1(44,60)            <= s_out1(45,60);
	s_locks_lower_in(44,60) <= s_locks_lower_out(45,60);

		normal_cell_45_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,1),
			fetch              => s_fetch(45,1),
			data_in            => s_data_in(45,1),
			data_out           => s_data_out(45,1),
			out1               => s_out1(45,1),
			out2               => s_out2(45,1),
			lock_lower_row_out => s_locks_lower_out(45,1),
			lock_lower_row_in  => s_locks_lower_in(45,1),
			in1                => s_in1(45,1),
			in2                => s_in2(45,1),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(1)
		);
	s_in1(45,1)            <= s_out1(46,1);
	s_in2(45,1)            <= s_out2(46,2);
	s_locks_lower_in(45,1) <= s_locks_lower_out(46,1);

		normal_cell_45_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,2),
			fetch              => s_fetch(45,2),
			data_in            => s_data_in(45,2),
			data_out           => s_data_out(45,2),
			out1               => s_out1(45,2),
			out2               => s_out2(45,2),
			lock_lower_row_out => s_locks_lower_out(45,2),
			lock_lower_row_in  => s_locks_lower_in(45,2),
			in1                => s_in1(45,2),
			in2                => s_in2(45,2),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(2)
		);
	s_in1(45,2)            <= s_out1(46,2);
	s_in2(45,2)            <= s_out2(46,3);
	s_locks_lower_in(45,2) <= s_locks_lower_out(46,2);

		normal_cell_45_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,3),
			fetch              => s_fetch(45,3),
			data_in            => s_data_in(45,3),
			data_out           => s_data_out(45,3),
			out1               => s_out1(45,3),
			out2               => s_out2(45,3),
			lock_lower_row_out => s_locks_lower_out(45,3),
			lock_lower_row_in  => s_locks_lower_in(45,3),
			in1                => s_in1(45,3),
			in2                => s_in2(45,3),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(3)
		);
	s_in1(45,3)            <= s_out1(46,3);
	s_in2(45,3)            <= s_out2(46,4);
	s_locks_lower_in(45,3) <= s_locks_lower_out(46,3);

		normal_cell_45_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,4),
			fetch              => s_fetch(45,4),
			data_in            => s_data_in(45,4),
			data_out           => s_data_out(45,4),
			out1               => s_out1(45,4),
			out2               => s_out2(45,4),
			lock_lower_row_out => s_locks_lower_out(45,4),
			lock_lower_row_in  => s_locks_lower_in(45,4),
			in1                => s_in1(45,4),
			in2                => s_in2(45,4),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(4)
		);
	s_in1(45,4)            <= s_out1(46,4);
	s_in2(45,4)            <= s_out2(46,5);
	s_locks_lower_in(45,4) <= s_locks_lower_out(46,4);

		normal_cell_45_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,5),
			fetch              => s_fetch(45,5),
			data_in            => s_data_in(45,5),
			data_out           => s_data_out(45,5),
			out1               => s_out1(45,5),
			out2               => s_out2(45,5),
			lock_lower_row_out => s_locks_lower_out(45,5),
			lock_lower_row_in  => s_locks_lower_in(45,5),
			in1                => s_in1(45,5),
			in2                => s_in2(45,5),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(5)
		);
	s_in1(45,5)            <= s_out1(46,5);
	s_in2(45,5)            <= s_out2(46,6);
	s_locks_lower_in(45,5) <= s_locks_lower_out(46,5);

		normal_cell_45_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,6),
			fetch              => s_fetch(45,6),
			data_in            => s_data_in(45,6),
			data_out           => s_data_out(45,6),
			out1               => s_out1(45,6),
			out2               => s_out2(45,6),
			lock_lower_row_out => s_locks_lower_out(45,6),
			lock_lower_row_in  => s_locks_lower_in(45,6),
			in1                => s_in1(45,6),
			in2                => s_in2(45,6),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(6)
		);
	s_in1(45,6)            <= s_out1(46,6);
	s_in2(45,6)            <= s_out2(46,7);
	s_locks_lower_in(45,6) <= s_locks_lower_out(46,6);

		normal_cell_45_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,7),
			fetch              => s_fetch(45,7),
			data_in            => s_data_in(45,7),
			data_out           => s_data_out(45,7),
			out1               => s_out1(45,7),
			out2               => s_out2(45,7),
			lock_lower_row_out => s_locks_lower_out(45,7),
			lock_lower_row_in  => s_locks_lower_in(45,7),
			in1                => s_in1(45,7),
			in2                => s_in2(45,7),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(7)
		);
	s_in1(45,7)            <= s_out1(46,7);
	s_in2(45,7)            <= s_out2(46,8);
	s_locks_lower_in(45,7) <= s_locks_lower_out(46,7);

		normal_cell_45_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,8),
			fetch              => s_fetch(45,8),
			data_in            => s_data_in(45,8),
			data_out           => s_data_out(45,8),
			out1               => s_out1(45,8),
			out2               => s_out2(45,8),
			lock_lower_row_out => s_locks_lower_out(45,8),
			lock_lower_row_in  => s_locks_lower_in(45,8),
			in1                => s_in1(45,8),
			in2                => s_in2(45,8),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(8)
		);
	s_in1(45,8)            <= s_out1(46,8);
	s_in2(45,8)            <= s_out2(46,9);
	s_locks_lower_in(45,8) <= s_locks_lower_out(46,8);

		normal_cell_45_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,9),
			fetch              => s_fetch(45,9),
			data_in            => s_data_in(45,9),
			data_out           => s_data_out(45,9),
			out1               => s_out1(45,9),
			out2               => s_out2(45,9),
			lock_lower_row_out => s_locks_lower_out(45,9),
			lock_lower_row_in  => s_locks_lower_in(45,9),
			in1                => s_in1(45,9),
			in2                => s_in2(45,9),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(9)
		);
	s_in1(45,9)            <= s_out1(46,9);
	s_in2(45,9)            <= s_out2(46,10);
	s_locks_lower_in(45,9) <= s_locks_lower_out(46,9);

		normal_cell_45_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,10),
			fetch              => s_fetch(45,10),
			data_in            => s_data_in(45,10),
			data_out           => s_data_out(45,10),
			out1               => s_out1(45,10),
			out2               => s_out2(45,10),
			lock_lower_row_out => s_locks_lower_out(45,10),
			lock_lower_row_in  => s_locks_lower_in(45,10),
			in1                => s_in1(45,10),
			in2                => s_in2(45,10),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(10)
		);
	s_in1(45,10)            <= s_out1(46,10);
	s_in2(45,10)            <= s_out2(46,11);
	s_locks_lower_in(45,10) <= s_locks_lower_out(46,10);

		normal_cell_45_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,11),
			fetch              => s_fetch(45,11),
			data_in            => s_data_in(45,11),
			data_out           => s_data_out(45,11),
			out1               => s_out1(45,11),
			out2               => s_out2(45,11),
			lock_lower_row_out => s_locks_lower_out(45,11),
			lock_lower_row_in  => s_locks_lower_in(45,11),
			in1                => s_in1(45,11),
			in2                => s_in2(45,11),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(11)
		);
	s_in1(45,11)            <= s_out1(46,11);
	s_in2(45,11)            <= s_out2(46,12);
	s_locks_lower_in(45,11) <= s_locks_lower_out(46,11);

		normal_cell_45_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,12),
			fetch              => s_fetch(45,12),
			data_in            => s_data_in(45,12),
			data_out           => s_data_out(45,12),
			out1               => s_out1(45,12),
			out2               => s_out2(45,12),
			lock_lower_row_out => s_locks_lower_out(45,12),
			lock_lower_row_in  => s_locks_lower_in(45,12),
			in1                => s_in1(45,12),
			in2                => s_in2(45,12),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(12)
		);
	s_in1(45,12)            <= s_out1(46,12);
	s_in2(45,12)            <= s_out2(46,13);
	s_locks_lower_in(45,12) <= s_locks_lower_out(46,12);

		normal_cell_45_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,13),
			fetch              => s_fetch(45,13),
			data_in            => s_data_in(45,13),
			data_out           => s_data_out(45,13),
			out1               => s_out1(45,13),
			out2               => s_out2(45,13),
			lock_lower_row_out => s_locks_lower_out(45,13),
			lock_lower_row_in  => s_locks_lower_in(45,13),
			in1                => s_in1(45,13),
			in2                => s_in2(45,13),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(13)
		);
	s_in1(45,13)            <= s_out1(46,13);
	s_in2(45,13)            <= s_out2(46,14);
	s_locks_lower_in(45,13) <= s_locks_lower_out(46,13);

		normal_cell_45_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,14),
			fetch              => s_fetch(45,14),
			data_in            => s_data_in(45,14),
			data_out           => s_data_out(45,14),
			out1               => s_out1(45,14),
			out2               => s_out2(45,14),
			lock_lower_row_out => s_locks_lower_out(45,14),
			lock_lower_row_in  => s_locks_lower_in(45,14),
			in1                => s_in1(45,14),
			in2                => s_in2(45,14),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(14)
		);
	s_in1(45,14)            <= s_out1(46,14);
	s_in2(45,14)            <= s_out2(46,15);
	s_locks_lower_in(45,14) <= s_locks_lower_out(46,14);

		normal_cell_45_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,15),
			fetch              => s_fetch(45,15),
			data_in            => s_data_in(45,15),
			data_out           => s_data_out(45,15),
			out1               => s_out1(45,15),
			out2               => s_out2(45,15),
			lock_lower_row_out => s_locks_lower_out(45,15),
			lock_lower_row_in  => s_locks_lower_in(45,15),
			in1                => s_in1(45,15),
			in2                => s_in2(45,15),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(15)
		);
	s_in1(45,15)            <= s_out1(46,15);
	s_in2(45,15)            <= s_out2(46,16);
	s_locks_lower_in(45,15) <= s_locks_lower_out(46,15);

		normal_cell_45_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,16),
			fetch              => s_fetch(45,16),
			data_in            => s_data_in(45,16),
			data_out           => s_data_out(45,16),
			out1               => s_out1(45,16),
			out2               => s_out2(45,16),
			lock_lower_row_out => s_locks_lower_out(45,16),
			lock_lower_row_in  => s_locks_lower_in(45,16),
			in1                => s_in1(45,16),
			in2                => s_in2(45,16),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(16)
		);
	s_in1(45,16)            <= s_out1(46,16);
	s_in2(45,16)            <= s_out2(46,17);
	s_locks_lower_in(45,16) <= s_locks_lower_out(46,16);

		normal_cell_45_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,17),
			fetch              => s_fetch(45,17),
			data_in            => s_data_in(45,17),
			data_out           => s_data_out(45,17),
			out1               => s_out1(45,17),
			out2               => s_out2(45,17),
			lock_lower_row_out => s_locks_lower_out(45,17),
			lock_lower_row_in  => s_locks_lower_in(45,17),
			in1                => s_in1(45,17),
			in2                => s_in2(45,17),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(17)
		);
	s_in1(45,17)            <= s_out1(46,17);
	s_in2(45,17)            <= s_out2(46,18);
	s_locks_lower_in(45,17) <= s_locks_lower_out(46,17);

		normal_cell_45_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,18),
			fetch              => s_fetch(45,18),
			data_in            => s_data_in(45,18),
			data_out           => s_data_out(45,18),
			out1               => s_out1(45,18),
			out2               => s_out2(45,18),
			lock_lower_row_out => s_locks_lower_out(45,18),
			lock_lower_row_in  => s_locks_lower_in(45,18),
			in1                => s_in1(45,18),
			in2                => s_in2(45,18),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(18)
		);
	s_in1(45,18)            <= s_out1(46,18);
	s_in2(45,18)            <= s_out2(46,19);
	s_locks_lower_in(45,18) <= s_locks_lower_out(46,18);

		normal_cell_45_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,19),
			fetch              => s_fetch(45,19),
			data_in            => s_data_in(45,19),
			data_out           => s_data_out(45,19),
			out1               => s_out1(45,19),
			out2               => s_out2(45,19),
			lock_lower_row_out => s_locks_lower_out(45,19),
			lock_lower_row_in  => s_locks_lower_in(45,19),
			in1                => s_in1(45,19),
			in2                => s_in2(45,19),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(19)
		);
	s_in1(45,19)            <= s_out1(46,19);
	s_in2(45,19)            <= s_out2(46,20);
	s_locks_lower_in(45,19) <= s_locks_lower_out(46,19);

		normal_cell_45_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,20),
			fetch              => s_fetch(45,20),
			data_in            => s_data_in(45,20),
			data_out           => s_data_out(45,20),
			out1               => s_out1(45,20),
			out2               => s_out2(45,20),
			lock_lower_row_out => s_locks_lower_out(45,20),
			lock_lower_row_in  => s_locks_lower_in(45,20),
			in1                => s_in1(45,20),
			in2                => s_in2(45,20),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(20)
		);
	s_in1(45,20)            <= s_out1(46,20);
	s_in2(45,20)            <= s_out2(46,21);
	s_locks_lower_in(45,20) <= s_locks_lower_out(46,20);

		normal_cell_45_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,21),
			fetch              => s_fetch(45,21),
			data_in            => s_data_in(45,21),
			data_out           => s_data_out(45,21),
			out1               => s_out1(45,21),
			out2               => s_out2(45,21),
			lock_lower_row_out => s_locks_lower_out(45,21),
			lock_lower_row_in  => s_locks_lower_in(45,21),
			in1                => s_in1(45,21),
			in2                => s_in2(45,21),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(21)
		);
	s_in1(45,21)            <= s_out1(46,21);
	s_in2(45,21)            <= s_out2(46,22);
	s_locks_lower_in(45,21) <= s_locks_lower_out(46,21);

		normal_cell_45_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,22),
			fetch              => s_fetch(45,22),
			data_in            => s_data_in(45,22),
			data_out           => s_data_out(45,22),
			out1               => s_out1(45,22),
			out2               => s_out2(45,22),
			lock_lower_row_out => s_locks_lower_out(45,22),
			lock_lower_row_in  => s_locks_lower_in(45,22),
			in1                => s_in1(45,22),
			in2                => s_in2(45,22),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(22)
		);
	s_in1(45,22)            <= s_out1(46,22);
	s_in2(45,22)            <= s_out2(46,23);
	s_locks_lower_in(45,22) <= s_locks_lower_out(46,22);

		normal_cell_45_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,23),
			fetch              => s_fetch(45,23),
			data_in            => s_data_in(45,23),
			data_out           => s_data_out(45,23),
			out1               => s_out1(45,23),
			out2               => s_out2(45,23),
			lock_lower_row_out => s_locks_lower_out(45,23),
			lock_lower_row_in  => s_locks_lower_in(45,23),
			in1                => s_in1(45,23),
			in2                => s_in2(45,23),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(23)
		);
	s_in1(45,23)            <= s_out1(46,23);
	s_in2(45,23)            <= s_out2(46,24);
	s_locks_lower_in(45,23) <= s_locks_lower_out(46,23);

		normal_cell_45_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,24),
			fetch              => s_fetch(45,24),
			data_in            => s_data_in(45,24),
			data_out           => s_data_out(45,24),
			out1               => s_out1(45,24),
			out2               => s_out2(45,24),
			lock_lower_row_out => s_locks_lower_out(45,24),
			lock_lower_row_in  => s_locks_lower_in(45,24),
			in1                => s_in1(45,24),
			in2                => s_in2(45,24),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(24)
		);
	s_in1(45,24)            <= s_out1(46,24);
	s_in2(45,24)            <= s_out2(46,25);
	s_locks_lower_in(45,24) <= s_locks_lower_out(46,24);

		normal_cell_45_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,25),
			fetch              => s_fetch(45,25),
			data_in            => s_data_in(45,25),
			data_out           => s_data_out(45,25),
			out1               => s_out1(45,25),
			out2               => s_out2(45,25),
			lock_lower_row_out => s_locks_lower_out(45,25),
			lock_lower_row_in  => s_locks_lower_in(45,25),
			in1                => s_in1(45,25),
			in2                => s_in2(45,25),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(25)
		);
	s_in1(45,25)            <= s_out1(46,25);
	s_in2(45,25)            <= s_out2(46,26);
	s_locks_lower_in(45,25) <= s_locks_lower_out(46,25);

		normal_cell_45_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,26),
			fetch              => s_fetch(45,26),
			data_in            => s_data_in(45,26),
			data_out           => s_data_out(45,26),
			out1               => s_out1(45,26),
			out2               => s_out2(45,26),
			lock_lower_row_out => s_locks_lower_out(45,26),
			lock_lower_row_in  => s_locks_lower_in(45,26),
			in1                => s_in1(45,26),
			in2                => s_in2(45,26),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(26)
		);
	s_in1(45,26)            <= s_out1(46,26);
	s_in2(45,26)            <= s_out2(46,27);
	s_locks_lower_in(45,26) <= s_locks_lower_out(46,26);

		normal_cell_45_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,27),
			fetch              => s_fetch(45,27),
			data_in            => s_data_in(45,27),
			data_out           => s_data_out(45,27),
			out1               => s_out1(45,27),
			out2               => s_out2(45,27),
			lock_lower_row_out => s_locks_lower_out(45,27),
			lock_lower_row_in  => s_locks_lower_in(45,27),
			in1                => s_in1(45,27),
			in2                => s_in2(45,27),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(27)
		);
	s_in1(45,27)            <= s_out1(46,27);
	s_in2(45,27)            <= s_out2(46,28);
	s_locks_lower_in(45,27) <= s_locks_lower_out(46,27);

		normal_cell_45_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,28),
			fetch              => s_fetch(45,28),
			data_in            => s_data_in(45,28),
			data_out           => s_data_out(45,28),
			out1               => s_out1(45,28),
			out2               => s_out2(45,28),
			lock_lower_row_out => s_locks_lower_out(45,28),
			lock_lower_row_in  => s_locks_lower_in(45,28),
			in1                => s_in1(45,28),
			in2                => s_in2(45,28),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(28)
		);
	s_in1(45,28)            <= s_out1(46,28);
	s_in2(45,28)            <= s_out2(46,29);
	s_locks_lower_in(45,28) <= s_locks_lower_out(46,28);

		normal_cell_45_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,29),
			fetch              => s_fetch(45,29),
			data_in            => s_data_in(45,29),
			data_out           => s_data_out(45,29),
			out1               => s_out1(45,29),
			out2               => s_out2(45,29),
			lock_lower_row_out => s_locks_lower_out(45,29),
			lock_lower_row_in  => s_locks_lower_in(45,29),
			in1                => s_in1(45,29),
			in2                => s_in2(45,29),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(29)
		);
	s_in1(45,29)            <= s_out1(46,29);
	s_in2(45,29)            <= s_out2(46,30);
	s_locks_lower_in(45,29) <= s_locks_lower_out(46,29);

		normal_cell_45_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,30),
			fetch              => s_fetch(45,30),
			data_in            => s_data_in(45,30),
			data_out           => s_data_out(45,30),
			out1               => s_out1(45,30),
			out2               => s_out2(45,30),
			lock_lower_row_out => s_locks_lower_out(45,30),
			lock_lower_row_in  => s_locks_lower_in(45,30),
			in1                => s_in1(45,30),
			in2                => s_in2(45,30),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(30)
		);
	s_in1(45,30)            <= s_out1(46,30);
	s_in2(45,30)            <= s_out2(46,31);
	s_locks_lower_in(45,30) <= s_locks_lower_out(46,30);

		normal_cell_45_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,31),
			fetch              => s_fetch(45,31),
			data_in            => s_data_in(45,31),
			data_out           => s_data_out(45,31),
			out1               => s_out1(45,31),
			out2               => s_out2(45,31),
			lock_lower_row_out => s_locks_lower_out(45,31),
			lock_lower_row_in  => s_locks_lower_in(45,31),
			in1                => s_in1(45,31),
			in2                => s_in2(45,31),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(31)
		);
	s_in1(45,31)            <= s_out1(46,31);
	s_in2(45,31)            <= s_out2(46,32);
	s_locks_lower_in(45,31) <= s_locks_lower_out(46,31);

		normal_cell_45_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,32),
			fetch              => s_fetch(45,32),
			data_in            => s_data_in(45,32),
			data_out           => s_data_out(45,32),
			out1               => s_out1(45,32),
			out2               => s_out2(45,32),
			lock_lower_row_out => s_locks_lower_out(45,32),
			lock_lower_row_in  => s_locks_lower_in(45,32),
			in1                => s_in1(45,32),
			in2                => s_in2(45,32),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(32)
		);
	s_in1(45,32)            <= s_out1(46,32);
	s_in2(45,32)            <= s_out2(46,33);
	s_locks_lower_in(45,32) <= s_locks_lower_out(46,32);

		normal_cell_45_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,33),
			fetch              => s_fetch(45,33),
			data_in            => s_data_in(45,33),
			data_out           => s_data_out(45,33),
			out1               => s_out1(45,33),
			out2               => s_out2(45,33),
			lock_lower_row_out => s_locks_lower_out(45,33),
			lock_lower_row_in  => s_locks_lower_in(45,33),
			in1                => s_in1(45,33),
			in2                => s_in2(45,33),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(33)
		);
	s_in1(45,33)            <= s_out1(46,33);
	s_in2(45,33)            <= s_out2(46,34);
	s_locks_lower_in(45,33) <= s_locks_lower_out(46,33);

		normal_cell_45_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,34),
			fetch              => s_fetch(45,34),
			data_in            => s_data_in(45,34),
			data_out           => s_data_out(45,34),
			out1               => s_out1(45,34),
			out2               => s_out2(45,34),
			lock_lower_row_out => s_locks_lower_out(45,34),
			lock_lower_row_in  => s_locks_lower_in(45,34),
			in1                => s_in1(45,34),
			in2                => s_in2(45,34),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(34)
		);
	s_in1(45,34)            <= s_out1(46,34);
	s_in2(45,34)            <= s_out2(46,35);
	s_locks_lower_in(45,34) <= s_locks_lower_out(46,34);

		normal_cell_45_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,35),
			fetch              => s_fetch(45,35),
			data_in            => s_data_in(45,35),
			data_out           => s_data_out(45,35),
			out1               => s_out1(45,35),
			out2               => s_out2(45,35),
			lock_lower_row_out => s_locks_lower_out(45,35),
			lock_lower_row_in  => s_locks_lower_in(45,35),
			in1                => s_in1(45,35),
			in2                => s_in2(45,35),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(35)
		);
	s_in1(45,35)            <= s_out1(46,35);
	s_in2(45,35)            <= s_out2(46,36);
	s_locks_lower_in(45,35) <= s_locks_lower_out(46,35);

		normal_cell_45_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,36),
			fetch              => s_fetch(45,36),
			data_in            => s_data_in(45,36),
			data_out           => s_data_out(45,36),
			out1               => s_out1(45,36),
			out2               => s_out2(45,36),
			lock_lower_row_out => s_locks_lower_out(45,36),
			lock_lower_row_in  => s_locks_lower_in(45,36),
			in1                => s_in1(45,36),
			in2                => s_in2(45,36),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(36)
		);
	s_in1(45,36)            <= s_out1(46,36);
	s_in2(45,36)            <= s_out2(46,37);
	s_locks_lower_in(45,36) <= s_locks_lower_out(46,36);

		normal_cell_45_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,37),
			fetch              => s_fetch(45,37),
			data_in            => s_data_in(45,37),
			data_out           => s_data_out(45,37),
			out1               => s_out1(45,37),
			out2               => s_out2(45,37),
			lock_lower_row_out => s_locks_lower_out(45,37),
			lock_lower_row_in  => s_locks_lower_in(45,37),
			in1                => s_in1(45,37),
			in2                => s_in2(45,37),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(37)
		);
	s_in1(45,37)            <= s_out1(46,37);
	s_in2(45,37)            <= s_out2(46,38);
	s_locks_lower_in(45,37) <= s_locks_lower_out(46,37);

		normal_cell_45_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,38),
			fetch              => s_fetch(45,38),
			data_in            => s_data_in(45,38),
			data_out           => s_data_out(45,38),
			out1               => s_out1(45,38),
			out2               => s_out2(45,38),
			lock_lower_row_out => s_locks_lower_out(45,38),
			lock_lower_row_in  => s_locks_lower_in(45,38),
			in1                => s_in1(45,38),
			in2                => s_in2(45,38),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(38)
		);
	s_in1(45,38)            <= s_out1(46,38);
	s_in2(45,38)            <= s_out2(46,39);
	s_locks_lower_in(45,38) <= s_locks_lower_out(46,38);

		normal_cell_45_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,39),
			fetch              => s_fetch(45,39),
			data_in            => s_data_in(45,39),
			data_out           => s_data_out(45,39),
			out1               => s_out1(45,39),
			out2               => s_out2(45,39),
			lock_lower_row_out => s_locks_lower_out(45,39),
			lock_lower_row_in  => s_locks_lower_in(45,39),
			in1                => s_in1(45,39),
			in2                => s_in2(45,39),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(39)
		);
	s_in1(45,39)            <= s_out1(46,39);
	s_in2(45,39)            <= s_out2(46,40);
	s_locks_lower_in(45,39) <= s_locks_lower_out(46,39);

		normal_cell_45_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,40),
			fetch              => s_fetch(45,40),
			data_in            => s_data_in(45,40),
			data_out           => s_data_out(45,40),
			out1               => s_out1(45,40),
			out2               => s_out2(45,40),
			lock_lower_row_out => s_locks_lower_out(45,40),
			lock_lower_row_in  => s_locks_lower_in(45,40),
			in1                => s_in1(45,40),
			in2                => s_in2(45,40),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(40)
		);
	s_in1(45,40)            <= s_out1(46,40);
	s_in2(45,40)            <= s_out2(46,41);
	s_locks_lower_in(45,40) <= s_locks_lower_out(46,40);

		normal_cell_45_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,41),
			fetch              => s_fetch(45,41),
			data_in            => s_data_in(45,41),
			data_out           => s_data_out(45,41),
			out1               => s_out1(45,41),
			out2               => s_out2(45,41),
			lock_lower_row_out => s_locks_lower_out(45,41),
			lock_lower_row_in  => s_locks_lower_in(45,41),
			in1                => s_in1(45,41),
			in2                => s_in2(45,41),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(41)
		);
	s_in1(45,41)            <= s_out1(46,41);
	s_in2(45,41)            <= s_out2(46,42);
	s_locks_lower_in(45,41) <= s_locks_lower_out(46,41);

		normal_cell_45_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,42),
			fetch              => s_fetch(45,42),
			data_in            => s_data_in(45,42),
			data_out           => s_data_out(45,42),
			out1               => s_out1(45,42),
			out2               => s_out2(45,42),
			lock_lower_row_out => s_locks_lower_out(45,42),
			lock_lower_row_in  => s_locks_lower_in(45,42),
			in1                => s_in1(45,42),
			in2                => s_in2(45,42),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(42)
		);
	s_in1(45,42)            <= s_out1(46,42);
	s_in2(45,42)            <= s_out2(46,43);
	s_locks_lower_in(45,42) <= s_locks_lower_out(46,42);

		normal_cell_45_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,43),
			fetch              => s_fetch(45,43),
			data_in            => s_data_in(45,43),
			data_out           => s_data_out(45,43),
			out1               => s_out1(45,43),
			out2               => s_out2(45,43),
			lock_lower_row_out => s_locks_lower_out(45,43),
			lock_lower_row_in  => s_locks_lower_in(45,43),
			in1                => s_in1(45,43),
			in2                => s_in2(45,43),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(43)
		);
	s_in1(45,43)            <= s_out1(46,43);
	s_in2(45,43)            <= s_out2(46,44);
	s_locks_lower_in(45,43) <= s_locks_lower_out(46,43);

		normal_cell_45_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,44),
			fetch              => s_fetch(45,44),
			data_in            => s_data_in(45,44),
			data_out           => s_data_out(45,44),
			out1               => s_out1(45,44),
			out2               => s_out2(45,44),
			lock_lower_row_out => s_locks_lower_out(45,44),
			lock_lower_row_in  => s_locks_lower_in(45,44),
			in1                => s_in1(45,44),
			in2                => s_in2(45,44),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(44)
		);
	s_in1(45,44)            <= s_out1(46,44);
	s_in2(45,44)            <= s_out2(46,45);
	s_locks_lower_in(45,44) <= s_locks_lower_out(46,44);

		normal_cell_45_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,45),
			fetch              => s_fetch(45,45),
			data_in            => s_data_in(45,45),
			data_out           => s_data_out(45,45),
			out1               => s_out1(45,45),
			out2               => s_out2(45,45),
			lock_lower_row_out => s_locks_lower_out(45,45),
			lock_lower_row_in  => s_locks_lower_in(45,45),
			in1                => s_in1(45,45),
			in2                => s_in2(45,45),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(45)
		);
	s_in1(45,45)            <= s_out1(46,45);
	s_in2(45,45)            <= s_out2(46,46);
	s_locks_lower_in(45,45) <= s_locks_lower_out(46,45);

		normal_cell_45_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,46),
			fetch              => s_fetch(45,46),
			data_in            => s_data_in(45,46),
			data_out           => s_data_out(45,46),
			out1               => s_out1(45,46),
			out2               => s_out2(45,46),
			lock_lower_row_out => s_locks_lower_out(45,46),
			lock_lower_row_in  => s_locks_lower_in(45,46),
			in1                => s_in1(45,46),
			in2                => s_in2(45,46),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(46)
		);
	s_in1(45,46)            <= s_out1(46,46);
	s_in2(45,46)            <= s_out2(46,47);
	s_locks_lower_in(45,46) <= s_locks_lower_out(46,46);

		normal_cell_45_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,47),
			fetch              => s_fetch(45,47),
			data_in            => s_data_in(45,47),
			data_out           => s_data_out(45,47),
			out1               => s_out1(45,47),
			out2               => s_out2(45,47),
			lock_lower_row_out => s_locks_lower_out(45,47),
			lock_lower_row_in  => s_locks_lower_in(45,47),
			in1                => s_in1(45,47),
			in2                => s_in2(45,47),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(47)
		);
	s_in1(45,47)            <= s_out1(46,47);
	s_in2(45,47)            <= s_out2(46,48);
	s_locks_lower_in(45,47) <= s_locks_lower_out(46,47);

		normal_cell_45_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,48),
			fetch              => s_fetch(45,48),
			data_in            => s_data_in(45,48),
			data_out           => s_data_out(45,48),
			out1               => s_out1(45,48),
			out2               => s_out2(45,48),
			lock_lower_row_out => s_locks_lower_out(45,48),
			lock_lower_row_in  => s_locks_lower_in(45,48),
			in1                => s_in1(45,48),
			in2                => s_in2(45,48),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(48)
		);
	s_in1(45,48)            <= s_out1(46,48);
	s_in2(45,48)            <= s_out2(46,49);
	s_locks_lower_in(45,48) <= s_locks_lower_out(46,48);

		normal_cell_45_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,49),
			fetch              => s_fetch(45,49),
			data_in            => s_data_in(45,49),
			data_out           => s_data_out(45,49),
			out1               => s_out1(45,49),
			out2               => s_out2(45,49),
			lock_lower_row_out => s_locks_lower_out(45,49),
			lock_lower_row_in  => s_locks_lower_in(45,49),
			in1                => s_in1(45,49),
			in2                => s_in2(45,49),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(49)
		);
	s_in1(45,49)            <= s_out1(46,49);
	s_in2(45,49)            <= s_out2(46,50);
	s_locks_lower_in(45,49) <= s_locks_lower_out(46,49);

		normal_cell_45_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,50),
			fetch              => s_fetch(45,50),
			data_in            => s_data_in(45,50),
			data_out           => s_data_out(45,50),
			out1               => s_out1(45,50),
			out2               => s_out2(45,50),
			lock_lower_row_out => s_locks_lower_out(45,50),
			lock_lower_row_in  => s_locks_lower_in(45,50),
			in1                => s_in1(45,50),
			in2                => s_in2(45,50),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(50)
		);
	s_in1(45,50)            <= s_out1(46,50);
	s_in2(45,50)            <= s_out2(46,51);
	s_locks_lower_in(45,50) <= s_locks_lower_out(46,50);

		normal_cell_45_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,51),
			fetch              => s_fetch(45,51),
			data_in            => s_data_in(45,51),
			data_out           => s_data_out(45,51),
			out1               => s_out1(45,51),
			out2               => s_out2(45,51),
			lock_lower_row_out => s_locks_lower_out(45,51),
			lock_lower_row_in  => s_locks_lower_in(45,51),
			in1                => s_in1(45,51),
			in2                => s_in2(45,51),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(51)
		);
	s_in1(45,51)            <= s_out1(46,51);
	s_in2(45,51)            <= s_out2(46,52);
	s_locks_lower_in(45,51) <= s_locks_lower_out(46,51);

		normal_cell_45_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,52),
			fetch              => s_fetch(45,52),
			data_in            => s_data_in(45,52),
			data_out           => s_data_out(45,52),
			out1               => s_out1(45,52),
			out2               => s_out2(45,52),
			lock_lower_row_out => s_locks_lower_out(45,52),
			lock_lower_row_in  => s_locks_lower_in(45,52),
			in1                => s_in1(45,52),
			in2                => s_in2(45,52),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(52)
		);
	s_in1(45,52)            <= s_out1(46,52);
	s_in2(45,52)            <= s_out2(46,53);
	s_locks_lower_in(45,52) <= s_locks_lower_out(46,52);

		normal_cell_45_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,53),
			fetch              => s_fetch(45,53),
			data_in            => s_data_in(45,53),
			data_out           => s_data_out(45,53),
			out1               => s_out1(45,53),
			out2               => s_out2(45,53),
			lock_lower_row_out => s_locks_lower_out(45,53),
			lock_lower_row_in  => s_locks_lower_in(45,53),
			in1                => s_in1(45,53),
			in2                => s_in2(45,53),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(53)
		);
	s_in1(45,53)            <= s_out1(46,53);
	s_in2(45,53)            <= s_out2(46,54);
	s_locks_lower_in(45,53) <= s_locks_lower_out(46,53);

		normal_cell_45_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,54),
			fetch              => s_fetch(45,54),
			data_in            => s_data_in(45,54),
			data_out           => s_data_out(45,54),
			out1               => s_out1(45,54),
			out2               => s_out2(45,54),
			lock_lower_row_out => s_locks_lower_out(45,54),
			lock_lower_row_in  => s_locks_lower_in(45,54),
			in1                => s_in1(45,54),
			in2                => s_in2(45,54),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(54)
		);
	s_in1(45,54)            <= s_out1(46,54);
	s_in2(45,54)            <= s_out2(46,55);
	s_locks_lower_in(45,54) <= s_locks_lower_out(46,54);

		normal_cell_45_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,55),
			fetch              => s_fetch(45,55),
			data_in            => s_data_in(45,55),
			data_out           => s_data_out(45,55),
			out1               => s_out1(45,55),
			out2               => s_out2(45,55),
			lock_lower_row_out => s_locks_lower_out(45,55),
			lock_lower_row_in  => s_locks_lower_in(45,55),
			in1                => s_in1(45,55),
			in2                => s_in2(45,55),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(55)
		);
	s_in1(45,55)            <= s_out1(46,55);
	s_in2(45,55)            <= s_out2(46,56);
	s_locks_lower_in(45,55) <= s_locks_lower_out(46,55);

		normal_cell_45_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,56),
			fetch              => s_fetch(45,56),
			data_in            => s_data_in(45,56),
			data_out           => s_data_out(45,56),
			out1               => s_out1(45,56),
			out2               => s_out2(45,56),
			lock_lower_row_out => s_locks_lower_out(45,56),
			lock_lower_row_in  => s_locks_lower_in(45,56),
			in1                => s_in1(45,56),
			in2                => s_in2(45,56),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(56)
		);
	s_in1(45,56)            <= s_out1(46,56);
	s_in2(45,56)            <= s_out2(46,57);
	s_locks_lower_in(45,56) <= s_locks_lower_out(46,56);

		normal_cell_45_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,57),
			fetch              => s_fetch(45,57),
			data_in            => s_data_in(45,57),
			data_out           => s_data_out(45,57),
			out1               => s_out1(45,57),
			out2               => s_out2(45,57),
			lock_lower_row_out => s_locks_lower_out(45,57),
			lock_lower_row_in  => s_locks_lower_in(45,57),
			in1                => s_in1(45,57),
			in2                => s_in2(45,57),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(57)
		);
	s_in1(45,57)            <= s_out1(46,57);
	s_in2(45,57)            <= s_out2(46,58);
	s_locks_lower_in(45,57) <= s_locks_lower_out(46,57);

		normal_cell_45_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,58),
			fetch              => s_fetch(45,58),
			data_in            => s_data_in(45,58),
			data_out           => s_data_out(45,58),
			out1               => s_out1(45,58),
			out2               => s_out2(45,58),
			lock_lower_row_out => s_locks_lower_out(45,58),
			lock_lower_row_in  => s_locks_lower_in(45,58),
			in1                => s_in1(45,58),
			in2                => s_in2(45,58),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(58)
		);
	s_in1(45,58)            <= s_out1(46,58);
	s_in2(45,58)            <= s_out2(46,59);
	s_locks_lower_in(45,58) <= s_locks_lower_out(46,58);

		normal_cell_45_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,59),
			fetch              => s_fetch(45,59),
			data_in            => s_data_in(45,59),
			data_out           => s_data_out(45,59),
			out1               => s_out1(45,59),
			out2               => s_out2(45,59),
			lock_lower_row_out => s_locks_lower_out(45,59),
			lock_lower_row_in  => s_locks_lower_in(45,59),
			in1                => s_in1(45,59),
			in2                => s_in2(45,59),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(59)
		);
	s_in1(45,59)            <= s_out1(46,59);
	s_in2(45,59)            <= s_out2(46,60);
	s_locks_lower_in(45,59) <= s_locks_lower_out(46,59);

		last_col_cell_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(45,60),
			fetch              => s_fetch(45,60),
			data_in            => s_data_in(45,60),
			data_out           => s_data_out(45,60),
			out1               => s_out1(45,60),
			out2               => s_out2(45,60),
			lock_lower_row_out => s_locks_lower_out(45,60),
			lock_lower_row_in  => s_locks_lower_in(45,60),
			in1                => s_in1(45,60),
			in2                => (others => '0'),
			lock_row           => s_locks(45),
			piv_found          => s_piv_found,
			row_data           => s_row_data(45),
			col_data           => s_col_data(60)
		);
	s_in1(45,60)            <= s_out1(46,60);
	s_locks_lower_in(45,60) <= s_locks_lower_out(46,60);

		normal_cell_46_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,1),
			fetch              => s_fetch(46,1),
			data_in            => s_data_in(46,1),
			data_out           => s_data_out(46,1),
			out1               => s_out1(46,1),
			out2               => s_out2(46,1),
			lock_lower_row_out => s_locks_lower_out(46,1),
			lock_lower_row_in  => s_locks_lower_in(46,1),
			in1                => s_in1(46,1),
			in2                => s_in2(46,1),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(1)
		);
	s_in1(46,1)            <= s_out1(47,1);
	s_in2(46,1)            <= s_out2(47,2);
	s_locks_lower_in(46,1) <= s_locks_lower_out(47,1);

		normal_cell_46_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,2),
			fetch              => s_fetch(46,2),
			data_in            => s_data_in(46,2),
			data_out           => s_data_out(46,2),
			out1               => s_out1(46,2),
			out2               => s_out2(46,2),
			lock_lower_row_out => s_locks_lower_out(46,2),
			lock_lower_row_in  => s_locks_lower_in(46,2),
			in1                => s_in1(46,2),
			in2                => s_in2(46,2),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(2)
		);
	s_in1(46,2)            <= s_out1(47,2);
	s_in2(46,2)            <= s_out2(47,3);
	s_locks_lower_in(46,2) <= s_locks_lower_out(47,2);

		normal_cell_46_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,3),
			fetch              => s_fetch(46,3),
			data_in            => s_data_in(46,3),
			data_out           => s_data_out(46,3),
			out1               => s_out1(46,3),
			out2               => s_out2(46,3),
			lock_lower_row_out => s_locks_lower_out(46,3),
			lock_lower_row_in  => s_locks_lower_in(46,3),
			in1                => s_in1(46,3),
			in2                => s_in2(46,3),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(3)
		);
	s_in1(46,3)            <= s_out1(47,3);
	s_in2(46,3)            <= s_out2(47,4);
	s_locks_lower_in(46,3) <= s_locks_lower_out(47,3);

		normal_cell_46_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,4),
			fetch              => s_fetch(46,4),
			data_in            => s_data_in(46,4),
			data_out           => s_data_out(46,4),
			out1               => s_out1(46,4),
			out2               => s_out2(46,4),
			lock_lower_row_out => s_locks_lower_out(46,4),
			lock_lower_row_in  => s_locks_lower_in(46,4),
			in1                => s_in1(46,4),
			in2                => s_in2(46,4),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(4)
		);
	s_in1(46,4)            <= s_out1(47,4);
	s_in2(46,4)            <= s_out2(47,5);
	s_locks_lower_in(46,4) <= s_locks_lower_out(47,4);

		normal_cell_46_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,5),
			fetch              => s_fetch(46,5),
			data_in            => s_data_in(46,5),
			data_out           => s_data_out(46,5),
			out1               => s_out1(46,5),
			out2               => s_out2(46,5),
			lock_lower_row_out => s_locks_lower_out(46,5),
			lock_lower_row_in  => s_locks_lower_in(46,5),
			in1                => s_in1(46,5),
			in2                => s_in2(46,5),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(5)
		);
	s_in1(46,5)            <= s_out1(47,5);
	s_in2(46,5)            <= s_out2(47,6);
	s_locks_lower_in(46,5) <= s_locks_lower_out(47,5);

		normal_cell_46_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,6),
			fetch              => s_fetch(46,6),
			data_in            => s_data_in(46,6),
			data_out           => s_data_out(46,6),
			out1               => s_out1(46,6),
			out2               => s_out2(46,6),
			lock_lower_row_out => s_locks_lower_out(46,6),
			lock_lower_row_in  => s_locks_lower_in(46,6),
			in1                => s_in1(46,6),
			in2                => s_in2(46,6),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(6)
		);
	s_in1(46,6)            <= s_out1(47,6);
	s_in2(46,6)            <= s_out2(47,7);
	s_locks_lower_in(46,6) <= s_locks_lower_out(47,6);

		normal_cell_46_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,7),
			fetch              => s_fetch(46,7),
			data_in            => s_data_in(46,7),
			data_out           => s_data_out(46,7),
			out1               => s_out1(46,7),
			out2               => s_out2(46,7),
			lock_lower_row_out => s_locks_lower_out(46,7),
			lock_lower_row_in  => s_locks_lower_in(46,7),
			in1                => s_in1(46,7),
			in2                => s_in2(46,7),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(7)
		);
	s_in1(46,7)            <= s_out1(47,7);
	s_in2(46,7)            <= s_out2(47,8);
	s_locks_lower_in(46,7) <= s_locks_lower_out(47,7);

		normal_cell_46_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,8),
			fetch              => s_fetch(46,8),
			data_in            => s_data_in(46,8),
			data_out           => s_data_out(46,8),
			out1               => s_out1(46,8),
			out2               => s_out2(46,8),
			lock_lower_row_out => s_locks_lower_out(46,8),
			lock_lower_row_in  => s_locks_lower_in(46,8),
			in1                => s_in1(46,8),
			in2                => s_in2(46,8),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(8)
		);
	s_in1(46,8)            <= s_out1(47,8);
	s_in2(46,8)            <= s_out2(47,9);
	s_locks_lower_in(46,8) <= s_locks_lower_out(47,8);

		normal_cell_46_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,9),
			fetch              => s_fetch(46,9),
			data_in            => s_data_in(46,9),
			data_out           => s_data_out(46,9),
			out1               => s_out1(46,9),
			out2               => s_out2(46,9),
			lock_lower_row_out => s_locks_lower_out(46,9),
			lock_lower_row_in  => s_locks_lower_in(46,9),
			in1                => s_in1(46,9),
			in2                => s_in2(46,9),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(9)
		);
	s_in1(46,9)            <= s_out1(47,9);
	s_in2(46,9)            <= s_out2(47,10);
	s_locks_lower_in(46,9) <= s_locks_lower_out(47,9);

		normal_cell_46_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,10),
			fetch              => s_fetch(46,10),
			data_in            => s_data_in(46,10),
			data_out           => s_data_out(46,10),
			out1               => s_out1(46,10),
			out2               => s_out2(46,10),
			lock_lower_row_out => s_locks_lower_out(46,10),
			lock_lower_row_in  => s_locks_lower_in(46,10),
			in1                => s_in1(46,10),
			in2                => s_in2(46,10),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(10)
		);
	s_in1(46,10)            <= s_out1(47,10);
	s_in2(46,10)            <= s_out2(47,11);
	s_locks_lower_in(46,10) <= s_locks_lower_out(47,10);

		normal_cell_46_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,11),
			fetch              => s_fetch(46,11),
			data_in            => s_data_in(46,11),
			data_out           => s_data_out(46,11),
			out1               => s_out1(46,11),
			out2               => s_out2(46,11),
			lock_lower_row_out => s_locks_lower_out(46,11),
			lock_lower_row_in  => s_locks_lower_in(46,11),
			in1                => s_in1(46,11),
			in2                => s_in2(46,11),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(11)
		);
	s_in1(46,11)            <= s_out1(47,11);
	s_in2(46,11)            <= s_out2(47,12);
	s_locks_lower_in(46,11) <= s_locks_lower_out(47,11);

		normal_cell_46_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,12),
			fetch              => s_fetch(46,12),
			data_in            => s_data_in(46,12),
			data_out           => s_data_out(46,12),
			out1               => s_out1(46,12),
			out2               => s_out2(46,12),
			lock_lower_row_out => s_locks_lower_out(46,12),
			lock_lower_row_in  => s_locks_lower_in(46,12),
			in1                => s_in1(46,12),
			in2                => s_in2(46,12),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(12)
		);
	s_in1(46,12)            <= s_out1(47,12);
	s_in2(46,12)            <= s_out2(47,13);
	s_locks_lower_in(46,12) <= s_locks_lower_out(47,12);

		normal_cell_46_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,13),
			fetch              => s_fetch(46,13),
			data_in            => s_data_in(46,13),
			data_out           => s_data_out(46,13),
			out1               => s_out1(46,13),
			out2               => s_out2(46,13),
			lock_lower_row_out => s_locks_lower_out(46,13),
			lock_lower_row_in  => s_locks_lower_in(46,13),
			in1                => s_in1(46,13),
			in2                => s_in2(46,13),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(13)
		);
	s_in1(46,13)            <= s_out1(47,13);
	s_in2(46,13)            <= s_out2(47,14);
	s_locks_lower_in(46,13) <= s_locks_lower_out(47,13);

		normal_cell_46_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,14),
			fetch              => s_fetch(46,14),
			data_in            => s_data_in(46,14),
			data_out           => s_data_out(46,14),
			out1               => s_out1(46,14),
			out2               => s_out2(46,14),
			lock_lower_row_out => s_locks_lower_out(46,14),
			lock_lower_row_in  => s_locks_lower_in(46,14),
			in1                => s_in1(46,14),
			in2                => s_in2(46,14),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(14)
		);
	s_in1(46,14)            <= s_out1(47,14);
	s_in2(46,14)            <= s_out2(47,15);
	s_locks_lower_in(46,14) <= s_locks_lower_out(47,14);

		normal_cell_46_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,15),
			fetch              => s_fetch(46,15),
			data_in            => s_data_in(46,15),
			data_out           => s_data_out(46,15),
			out1               => s_out1(46,15),
			out2               => s_out2(46,15),
			lock_lower_row_out => s_locks_lower_out(46,15),
			lock_lower_row_in  => s_locks_lower_in(46,15),
			in1                => s_in1(46,15),
			in2                => s_in2(46,15),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(15)
		);
	s_in1(46,15)            <= s_out1(47,15);
	s_in2(46,15)            <= s_out2(47,16);
	s_locks_lower_in(46,15) <= s_locks_lower_out(47,15);

		normal_cell_46_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,16),
			fetch              => s_fetch(46,16),
			data_in            => s_data_in(46,16),
			data_out           => s_data_out(46,16),
			out1               => s_out1(46,16),
			out2               => s_out2(46,16),
			lock_lower_row_out => s_locks_lower_out(46,16),
			lock_lower_row_in  => s_locks_lower_in(46,16),
			in1                => s_in1(46,16),
			in2                => s_in2(46,16),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(16)
		);
	s_in1(46,16)            <= s_out1(47,16);
	s_in2(46,16)            <= s_out2(47,17);
	s_locks_lower_in(46,16) <= s_locks_lower_out(47,16);

		normal_cell_46_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,17),
			fetch              => s_fetch(46,17),
			data_in            => s_data_in(46,17),
			data_out           => s_data_out(46,17),
			out1               => s_out1(46,17),
			out2               => s_out2(46,17),
			lock_lower_row_out => s_locks_lower_out(46,17),
			lock_lower_row_in  => s_locks_lower_in(46,17),
			in1                => s_in1(46,17),
			in2                => s_in2(46,17),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(17)
		);
	s_in1(46,17)            <= s_out1(47,17);
	s_in2(46,17)            <= s_out2(47,18);
	s_locks_lower_in(46,17) <= s_locks_lower_out(47,17);

		normal_cell_46_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,18),
			fetch              => s_fetch(46,18),
			data_in            => s_data_in(46,18),
			data_out           => s_data_out(46,18),
			out1               => s_out1(46,18),
			out2               => s_out2(46,18),
			lock_lower_row_out => s_locks_lower_out(46,18),
			lock_lower_row_in  => s_locks_lower_in(46,18),
			in1                => s_in1(46,18),
			in2                => s_in2(46,18),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(18)
		);
	s_in1(46,18)            <= s_out1(47,18);
	s_in2(46,18)            <= s_out2(47,19);
	s_locks_lower_in(46,18) <= s_locks_lower_out(47,18);

		normal_cell_46_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,19),
			fetch              => s_fetch(46,19),
			data_in            => s_data_in(46,19),
			data_out           => s_data_out(46,19),
			out1               => s_out1(46,19),
			out2               => s_out2(46,19),
			lock_lower_row_out => s_locks_lower_out(46,19),
			lock_lower_row_in  => s_locks_lower_in(46,19),
			in1                => s_in1(46,19),
			in2                => s_in2(46,19),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(19)
		);
	s_in1(46,19)            <= s_out1(47,19);
	s_in2(46,19)            <= s_out2(47,20);
	s_locks_lower_in(46,19) <= s_locks_lower_out(47,19);

		normal_cell_46_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,20),
			fetch              => s_fetch(46,20),
			data_in            => s_data_in(46,20),
			data_out           => s_data_out(46,20),
			out1               => s_out1(46,20),
			out2               => s_out2(46,20),
			lock_lower_row_out => s_locks_lower_out(46,20),
			lock_lower_row_in  => s_locks_lower_in(46,20),
			in1                => s_in1(46,20),
			in2                => s_in2(46,20),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(20)
		);
	s_in1(46,20)            <= s_out1(47,20);
	s_in2(46,20)            <= s_out2(47,21);
	s_locks_lower_in(46,20) <= s_locks_lower_out(47,20);

		normal_cell_46_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,21),
			fetch              => s_fetch(46,21),
			data_in            => s_data_in(46,21),
			data_out           => s_data_out(46,21),
			out1               => s_out1(46,21),
			out2               => s_out2(46,21),
			lock_lower_row_out => s_locks_lower_out(46,21),
			lock_lower_row_in  => s_locks_lower_in(46,21),
			in1                => s_in1(46,21),
			in2                => s_in2(46,21),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(21)
		);
	s_in1(46,21)            <= s_out1(47,21);
	s_in2(46,21)            <= s_out2(47,22);
	s_locks_lower_in(46,21) <= s_locks_lower_out(47,21);

		normal_cell_46_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,22),
			fetch              => s_fetch(46,22),
			data_in            => s_data_in(46,22),
			data_out           => s_data_out(46,22),
			out1               => s_out1(46,22),
			out2               => s_out2(46,22),
			lock_lower_row_out => s_locks_lower_out(46,22),
			lock_lower_row_in  => s_locks_lower_in(46,22),
			in1                => s_in1(46,22),
			in2                => s_in2(46,22),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(22)
		);
	s_in1(46,22)            <= s_out1(47,22);
	s_in2(46,22)            <= s_out2(47,23);
	s_locks_lower_in(46,22) <= s_locks_lower_out(47,22);

		normal_cell_46_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,23),
			fetch              => s_fetch(46,23),
			data_in            => s_data_in(46,23),
			data_out           => s_data_out(46,23),
			out1               => s_out1(46,23),
			out2               => s_out2(46,23),
			lock_lower_row_out => s_locks_lower_out(46,23),
			lock_lower_row_in  => s_locks_lower_in(46,23),
			in1                => s_in1(46,23),
			in2                => s_in2(46,23),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(23)
		);
	s_in1(46,23)            <= s_out1(47,23);
	s_in2(46,23)            <= s_out2(47,24);
	s_locks_lower_in(46,23) <= s_locks_lower_out(47,23);

		normal_cell_46_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,24),
			fetch              => s_fetch(46,24),
			data_in            => s_data_in(46,24),
			data_out           => s_data_out(46,24),
			out1               => s_out1(46,24),
			out2               => s_out2(46,24),
			lock_lower_row_out => s_locks_lower_out(46,24),
			lock_lower_row_in  => s_locks_lower_in(46,24),
			in1                => s_in1(46,24),
			in2                => s_in2(46,24),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(24)
		);
	s_in1(46,24)            <= s_out1(47,24);
	s_in2(46,24)            <= s_out2(47,25);
	s_locks_lower_in(46,24) <= s_locks_lower_out(47,24);

		normal_cell_46_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,25),
			fetch              => s_fetch(46,25),
			data_in            => s_data_in(46,25),
			data_out           => s_data_out(46,25),
			out1               => s_out1(46,25),
			out2               => s_out2(46,25),
			lock_lower_row_out => s_locks_lower_out(46,25),
			lock_lower_row_in  => s_locks_lower_in(46,25),
			in1                => s_in1(46,25),
			in2                => s_in2(46,25),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(25)
		);
	s_in1(46,25)            <= s_out1(47,25);
	s_in2(46,25)            <= s_out2(47,26);
	s_locks_lower_in(46,25) <= s_locks_lower_out(47,25);

		normal_cell_46_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,26),
			fetch              => s_fetch(46,26),
			data_in            => s_data_in(46,26),
			data_out           => s_data_out(46,26),
			out1               => s_out1(46,26),
			out2               => s_out2(46,26),
			lock_lower_row_out => s_locks_lower_out(46,26),
			lock_lower_row_in  => s_locks_lower_in(46,26),
			in1                => s_in1(46,26),
			in2                => s_in2(46,26),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(26)
		);
	s_in1(46,26)            <= s_out1(47,26);
	s_in2(46,26)            <= s_out2(47,27);
	s_locks_lower_in(46,26) <= s_locks_lower_out(47,26);

		normal_cell_46_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,27),
			fetch              => s_fetch(46,27),
			data_in            => s_data_in(46,27),
			data_out           => s_data_out(46,27),
			out1               => s_out1(46,27),
			out2               => s_out2(46,27),
			lock_lower_row_out => s_locks_lower_out(46,27),
			lock_lower_row_in  => s_locks_lower_in(46,27),
			in1                => s_in1(46,27),
			in2                => s_in2(46,27),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(27)
		);
	s_in1(46,27)            <= s_out1(47,27);
	s_in2(46,27)            <= s_out2(47,28);
	s_locks_lower_in(46,27) <= s_locks_lower_out(47,27);

		normal_cell_46_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,28),
			fetch              => s_fetch(46,28),
			data_in            => s_data_in(46,28),
			data_out           => s_data_out(46,28),
			out1               => s_out1(46,28),
			out2               => s_out2(46,28),
			lock_lower_row_out => s_locks_lower_out(46,28),
			lock_lower_row_in  => s_locks_lower_in(46,28),
			in1                => s_in1(46,28),
			in2                => s_in2(46,28),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(28)
		);
	s_in1(46,28)            <= s_out1(47,28);
	s_in2(46,28)            <= s_out2(47,29);
	s_locks_lower_in(46,28) <= s_locks_lower_out(47,28);

		normal_cell_46_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,29),
			fetch              => s_fetch(46,29),
			data_in            => s_data_in(46,29),
			data_out           => s_data_out(46,29),
			out1               => s_out1(46,29),
			out2               => s_out2(46,29),
			lock_lower_row_out => s_locks_lower_out(46,29),
			lock_lower_row_in  => s_locks_lower_in(46,29),
			in1                => s_in1(46,29),
			in2                => s_in2(46,29),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(29)
		);
	s_in1(46,29)            <= s_out1(47,29);
	s_in2(46,29)            <= s_out2(47,30);
	s_locks_lower_in(46,29) <= s_locks_lower_out(47,29);

		normal_cell_46_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,30),
			fetch              => s_fetch(46,30),
			data_in            => s_data_in(46,30),
			data_out           => s_data_out(46,30),
			out1               => s_out1(46,30),
			out2               => s_out2(46,30),
			lock_lower_row_out => s_locks_lower_out(46,30),
			lock_lower_row_in  => s_locks_lower_in(46,30),
			in1                => s_in1(46,30),
			in2                => s_in2(46,30),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(30)
		);
	s_in1(46,30)            <= s_out1(47,30);
	s_in2(46,30)            <= s_out2(47,31);
	s_locks_lower_in(46,30) <= s_locks_lower_out(47,30);

		normal_cell_46_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,31),
			fetch              => s_fetch(46,31),
			data_in            => s_data_in(46,31),
			data_out           => s_data_out(46,31),
			out1               => s_out1(46,31),
			out2               => s_out2(46,31),
			lock_lower_row_out => s_locks_lower_out(46,31),
			lock_lower_row_in  => s_locks_lower_in(46,31),
			in1                => s_in1(46,31),
			in2                => s_in2(46,31),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(31)
		);
	s_in1(46,31)            <= s_out1(47,31);
	s_in2(46,31)            <= s_out2(47,32);
	s_locks_lower_in(46,31) <= s_locks_lower_out(47,31);

		normal_cell_46_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,32),
			fetch              => s_fetch(46,32),
			data_in            => s_data_in(46,32),
			data_out           => s_data_out(46,32),
			out1               => s_out1(46,32),
			out2               => s_out2(46,32),
			lock_lower_row_out => s_locks_lower_out(46,32),
			lock_lower_row_in  => s_locks_lower_in(46,32),
			in1                => s_in1(46,32),
			in2                => s_in2(46,32),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(32)
		);
	s_in1(46,32)            <= s_out1(47,32);
	s_in2(46,32)            <= s_out2(47,33);
	s_locks_lower_in(46,32) <= s_locks_lower_out(47,32);

		normal_cell_46_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,33),
			fetch              => s_fetch(46,33),
			data_in            => s_data_in(46,33),
			data_out           => s_data_out(46,33),
			out1               => s_out1(46,33),
			out2               => s_out2(46,33),
			lock_lower_row_out => s_locks_lower_out(46,33),
			lock_lower_row_in  => s_locks_lower_in(46,33),
			in1                => s_in1(46,33),
			in2                => s_in2(46,33),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(33)
		);
	s_in1(46,33)            <= s_out1(47,33);
	s_in2(46,33)            <= s_out2(47,34);
	s_locks_lower_in(46,33) <= s_locks_lower_out(47,33);

		normal_cell_46_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,34),
			fetch              => s_fetch(46,34),
			data_in            => s_data_in(46,34),
			data_out           => s_data_out(46,34),
			out1               => s_out1(46,34),
			out2               => s_out2(46,34),
			lock_lower_row_out => s_locks_lower_out(46,34),
			lock_lower_row_in  => s_locks_lower_in(46,34),
			in1                => s_in1(46,34),
			in2                => s_in2(46,34),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(34)
		);
	s_in1(46,34)            <= s_out1(47,34);
	s_in2(46,34)            <= s_out2(47,35);
	s_locks_lower_in(46,34) <= s_locks_lower_out(47,34);

		normal_cell_46_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,35),
			fetch              => s_fetch(46,35),
			data_in            => s_data_in(46,35),
			data_out           => s_data_out(46,35),
			out1               => s_out1(46,35),
			out2               => s_out2(46,35),
			lock_lower_row_out => s_locks_lower_out(46,35),
			lock_lower_row_in  => s_locks_lower_in(46,35),
			in1                => s_in1(46,35),
			in2                => s_in2(46,35),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(35)
		);
	s_in1(46,35)            <= s_out1(47,35);
	s_in2(46,35)            <= s_out2(47,36);
	s_locks_lower_in(46,35) <= s_locks_lower_out(47,35);

		normal_cell_46_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,36),
			fetch              => s_fetch(46,36),
			data_in            => s_data_in(46,36),
			data_out           => s_data_out(46,36),
			out1               => s_out1(46,36),
			out2               => s_out2(46,36),
			lock_lower_row_out => s_locks_lower_out(46,36),
			lock_lower_row_in  => s_locks_lower_in(46,36),
			in1                => s_in1(46,36),
			in2                => s_in2(46,36),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(36)
		);
	s_in1(46,36)            <= s_out1(47,36);
	s_in2(46,36)            <= s_out2(47,37);
	s_locks_lower_in(46,36) <= s_locks_lower_out(47,36);

		normal_cell_46_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,37),
			fetch              => s_fetch(46,37),
			data_in            => s_data_in(46,37),
			data_out           => s_data_out(46,37),
			out1               => s_out1(46,37),
			out2               => s_out2(46,37),
			lock_lower_row_out => s_locks_lower_out(46,37),
			lock_lower_row_in  => s_locks_lower_in(46,37),
			in1                => s_in1(46,37),
			in2                => s_in2(46,37),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(37)
		);
	s_in1(46,37)            <= s_out1(47,37);
	s_in2(46,37)            <= s_out2(47,38);
	s_locks_lower_in(46,37) <= s_locks_lower_out(47,37);

		normal_cell_46_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,38),
			fetch              => s_fetch(46,38),
			data_in            => s_data_in(46,38),
			data_out           => s_data_out(46,38),
			out1               => s_out1(46,38),
			out2               => s_out2(46,38),
			lock_lower_row_out => s_locks_lower_out(46,38),
			lock_lower_row_in  => s_locks_lower_in(46,38),
			in1                => s_in1(46,38),
			in2                => s_in2(46,38),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(38)
		);
	s_in1(46,38)            <= s_out1(47,38);
	s_in2(46,38)            <= s_out2(47,39);
	s_locks_lower_in(46,38) <= s_locks_lower_out(47,38);

		normal_cell_46_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,39),
			fetch              => s_fetch(46,39),
			data_in            => s_data_in(46,39),
			data_out           => s_data_out(46,39),
			out1               => s_out1(46,39),
			out2               => s_out2(46,39),
			lock_lower_row_out => s_locks_lower_out(46,39),
			lock_lower_row_in  => s_locks_lower_in(46,39),
			in1                => s_in1(46,39),
			in2                => s_in2(46,39),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(39)
		);
	s_in1(46,39)            <= s_out1(47,39);
	s_in2(46,39)            <= s_out2(47,40);
	s_locks_lower_in(46,39) <= s_locks_lower_out(47,39);

		normal_cell_46_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,40),
			fetch              => s_fetch(46,40),
			data_in            => s_data_in(46,40),
			data_out           => s_data_out(46,40),
			out1               => s_out1(46,40),
			out2               => s_out2(46,40),
			lock_lower_row_out => s_locks_lower_out(46,40),
			lock_lower_row_in  => s_locks_lower_in(46,40),
			in1                => s_in1(46,40),
			in2                => s_in2(46,40),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(40)
		);
	s_in1(46,40)            <= s_out1(47,40);
	s_in2(46,40)            <= s_out2(47,41);
	s_locks_lower_in(46,40) <= s_locks_lower_out(47,40);

		normal_cell_46_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,41),
			fetch              => s_fetch(46,41),
			data_in            => s_data_in(46,41),
			data_out           => s_data_out(46,41),
			out1               => s_out1(46,41),
			out2               => s_out2(46,41),
			lock_lower_row_out => s_locks_lower_out(46,41),
			lock_lower_row_in  => s_locks_lower_in(46,41),
			in1                => s_in1(46,41),
			in2                => s_in2(46,41),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(41)
		);
	s_in1(46,41)            <= s_out1(47,41);
	s_in2(46,41)            <= s_out2(47,42);
	s_locks_lower_in(46,41) <= s_locks_lower_out(47,41);

		normal_cell_46_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,42),
			fetch              => s_fetch(46,42),
			data_in            => s_data_in(46,42),
			data_out           => s_data_out(46,42),
			out1               => s_out1(46,42),
			out2               => s_out2(46,42),
			lock_lower_row_out => s_locks_lower_out(46,42),
			lock_lower_row_in  => s_locks_lower_in(46,42),
			in1                => s_in1(46,42),
			in2                => s_in2(46,42),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(42)
		);
	s_in1(46,42)            <= s_out1(47,42);
	s_in2(46,42)            <= s_out2(47,43);
	s_locks_lower_in(46,42) <= s_locks_lower_out(47,42);

		normal_cell_46_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,43),
			fetch              => s_fetch(46,43),
			data_in            => s_data_in(46,43),
			data_out           => s_data_out(46,43),
			out1               => s_out1(46,43),
			out2               => s_out2(46,43),
			lock_lower_row_out => s_locks_lower_out(46,43),
			lock_lower_row_in  => s_locks_lower_in(46,43),
			in1                => s_in1(46,43),
			in2                => s_in2(46,43),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(43)
		);
	s_in1(46,43)            <= s_out1(47,43);
	s_in2(46,43)            <= s_out2(47,44);
	s_locks_lower_in(46,43) <= s_locks_lower_out(47,43);

		normal_cell_46_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,44),
			fetch              => s_fetch(46,44),
			data_in            => s_data_in(46,44),
			data_out           => s_data_out(46,44),
			out1               => s_out1(46,44),
			out2               => s_out2(46,44),
			lock_lower_row_out => s_locks_lower_out(46,44),
			lock_lower_row_in  => s_locks_lower_in(46,44),
			in1                => s_in1(46,44),
			in2                => s_in2(46,44),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(44)
		);
	s_in1(46,44)            <= s_out1(47,44);
	s_in2(46,44)            <= s_out2(47,45);
	s_locks_lower_in(46,44) <= s_locks_lower_out(47,44);

		normal_cell_46_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,45),
			fetch              => s_fetch(46,45),
			data_in            => s_data_in(46,45),
			data_out           => s_data_out(46,45),
			out1               => s_out1(46,45),
			out2               => s_out2(46,45),
			lock_lower_row_out => s_locks_lower_out(46,45),
			lock_lower_row_in  => s_locks_lower_in(46,45),
			in1                => s_in1(46,45),
			in2                => s_in2(46,45),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(45)
		);
	s_in1(46,45)            <= s_out1(47,45);
	s_in2(46,45)            <= s_out2(47,46);
	s_locks_lower_in(46,45) <= s_locks_lower_out(47,45);

		normal_cell_46_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,46),
			fetch              => s_fetch(46,46),
			data_in            => s_data_in(46,46),
			data_out           => s_data_out(46,46),
			out1               => s_out1(46,46),
			out2               => s_out2(46,46),
			lock_lower_row_out => s_locks_lower_out(46,46),
			lock_lower_row_in  => s_locks_lower_in(46,46),
			in1                => s_in1(46,46),
			in2                => s_in2(46,46),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(46)
		);
	s_in1(46,46)            <= s_out1(47,46);
	s_in2(46,46)            <= s_out2(47,47);
	s_locks_lower_in(46,46) <= s_locks_lower_out(47,46);

		normal_cell_46_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,47),
			fetch              => s_fetch(46,47),
			data_in            => s_data_in(46,47),
			data_out           => s_data_out(46,47),
			out1               => s_out1(46,47),
			out2               => s_out2(46,47),
			lock_lower_row_out => s_locks_lower_out(46,47),
			lock_lower_row_in  => s_locks_lower_in(46,47),
			in1                => s_in1(46,47),
			in2                => s_in2(46,47),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(47)
		);
	s_in1(46,47)            <= s_out1(47,47);
	s_in2(46,47)            <= s_out2(47,48);
	s_locks_lower_in(46,47) <= s_locks_lower_out(47,47);

		normal_cell_46_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,48),
			fetch              => s_fetch(46,48),
			data_in            => s_data_in(46,48),
			data_out           => s_data_out(46,48),
			out1               => s_out1(46,48),
			out2               => s_out2(46,48),
			lock_lower_row_out => s_locks_lower_out(46,48),
			lock_lower_row_in  => s_locks_lower_in(46,48),
			in1                => s_in1(46,48),
			in2                => s_in2(46,48),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(48)
		);
	s_in1(46,48)            <= s_out1(47,48);
	s_in2(46,48)            <= s_out2(47,49);
	s_locks_lower_in(46,48) <= s_locks_lower_out(47,48);

		normal_cell_46_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,49),
			fetch              => s_fetch(46,49),
			data_in            => s_data_in(46,49),
			data_out           => s_data_out(46,49),
			out1               => s_out1(46,49),
			out2               => s_out2(46,49),
			lock_lower_row_out => s_locks_lower_out(46,49),
			lock_lower_row_in  => s_locks_lower_in(46,49),
			in1                => s_in1(46,49),
			in2                => s_in2(46,49),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(49)
		);
	s_in1(46,49)            <= s_out1(47,49);
	s_in2(46,49)            <= s_out2(47,50);
	s_locks_lower_in(46,49) <= s_locks_lower_out(47,49);

		normal_cell_46_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,50),
			fetch              => s_fetch(46,50),
			data_in            => s_data_in(46,50),
			data_out           => s_data_out(46,50),
			out1               => s_out1(46,50),
			out2               => s_out2(46,50),
			lock_lower_row_out => s_locks_lower_out(46,50),
			lock_lower_row_in  => s_locks_lower_in(46,50),
			in1                => s_in1(46,50),
			in2                => s_in2(46,50),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(50)
		);
	s_in1(46,50)            <= s_out1(47,50);
	s_in2(46,50)            <= s_out2(47,51);
	s_locks_lower_in(46,50) <= s_locks_lower_out(47,50);

		normal_cell_46_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,51),
			fetch              => s_fetch(46,51),
			data_in            => s_data_in(46,51),
			data_out           => s_data_out(46,51),
			out1               => s_out1(46,51),
			out2               => s_out2(46,51),
			lock_lower_row_out => s_locks_lower_out(46,51),
			lock_lower_row_in  => s_locks_lower_in(46,51),
			in1                => s_in1(46,51),
			in2                => s_in2(46,51),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(51)
		);
	s_in1(46,51)            <= s_out1(47,51);
	s_in2(46,51)            <= s_out2(47,52);
	s_locks_lower_in(46,51) <= s_locks_lower_out(47,51);

		normal_cell_46_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,52),
			fetch              => s_fetch(46,52),
			data_in            => s_data_in(46,52),
			data_out           => s_data_out(46,52),
			out1               => s_out1(46,52),
			out2               => s_out2(46,52),
			lock_lower_row_out => s_locks_lower_out(46,52),
			lock_lower_row_in  => s_locks_lower_in(46,52),
			in1                => s_in1(46,52),
			in2                => s_in2(46,52),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(52)
		);
	s_in1(46,52)            <= s_out1(47,52);
	s_in2(46,52)            <= s_out2(47,53);
	s_locks_lower_in(46,52) <= s_locks_lower_out(47,52);

		normal_cell_46_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,53),
			fetch              => s_fetch(46,53),
			data_in            => s_data_in(46,53),
			data_out           => s_data_out(46,53),
			out1               => s_out1(46,53),
			out2               => s_out2(46,53),
			lock_lower_row_out => s_locks_lower_out(46,53),
			lock_lower_row_in  => s_locks_lower_in(46,53),
			in1                => s_in1(46,53),
			in2                => s_in2(46,53),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(53)
		);
	s_in1(46,53)            <= s_out1(47,53);
	s_in2(46,53)            <= s_out2(47,54);
	s_locks_lower_in(46,53) <= s_locks_lower_out(47,53);

		normal_cell_46_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,54),
			fetch              => s_fetch(46,54),
			data_in            => s_data_in(46,54),
			data_out           => s_data_out(46,54),
			out1               => s_out1(46,54),
			out2               => s_out2(46,54),
			lock_lower_row_out => s_locks_lower_out(46,54),
			lock_lower_row_in  => s_locks_lower_in(46,54),
			in1                => s_in1(46,54),
			in2                => s_in2(46,54),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(54)
		);
	s_in1(46,54)            <= s_out1(47,54);
	s_in2(46,54)            <= s_out2(47,55);
	s_locks_lower_in(46,54) <= s_locks_lower_out(47,54);

		normal_cell_46_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,55),
			fetch              => s_fetch(46,55),
			data_in            => s_data_in(46,55),
			data_out           => s_data_out(46,55),
			out1               => s_out1(46,55),
			out2               => s_out2(46,55),
			lock_lower_row_out => s_locks_lower_out(46,55),
			lock_lower_row_in  => s_locks_lower_in(46,55),
			in1                => s_in1(46,55),
			in2                => s_in2(46,55),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(55)
		);
	s_in1(46,55)            <= s_out1(47,55);
	s_in2(46,55)            <= s_out2(47,56);
	s_locks_lower_in(46,55) <= s_locks_lower_out(47,55);

		normal_cell_46_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,56),
			fetch              => s_fetch(46,56),
			data_in            => s_data_in(46,56),
			data_out           => s_data_out(46,56),
			out1               => s_out1(46,56),
			out2               => s_out2(46,56),
			lock_lower_row_out => s_locks_lower_out(46,56),
			lock_lower_row_in  => s_locks_lower_in(46,56),
			in1                => s_in1(46,56),
			in2                => s_in2(46,56),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(56)
		);
	s_in1(46,56)            <= s_out1(47,56);
	s_in2(46,56)            <= s_out2(47,57);
	s_locks_lower_in(46,56) <= s_locks_lower_out(47,56);

		normal_cell_46_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,57),
			fetch              => s_fetch(46,57),
			data_in            => s_data_in(46,57),
			data_out           => s_data_out(46,57),
			out1               => s_out1(46,57),
			out2               => s_out2(46,57),
			lock_lower_row_out => s_locks_lower_out(46,57),
			lock_lower_row_in  => s_locks_lower_in(46,57),
			in1                => s_in1(46,57),
			in2                => s_in2(46,57),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(57)
		);
	s_in1(46,57)            <= s_out1(47,57);
	s_in2(46,57)            <= s_out2(47,58);
	s_locks_lower_in(46,57) <= s_locks_lower_out(47,57);

		normal_cell_46_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,58),
			fetch              => s_fetch(46,58),
			data_in            => s_data_in(46,58),
			data_out           => s_data_out(46,58),
			out1               => s_out1(46,58),
			out2               => s_out2(46,58),
			lock_lower_row_out => s_locks_lower_out(46,58),
			lock_lower_row_in  => s_locks_lower_in(46,58),
			in1                => s_in1(46,58),
			in2                => s_in2(46,58),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(58)
		);
	s_in1(46,58)            <= s_out1(47,58);
	s_in2(46,58)            <= s_out2(47,59);
	s_locks_lower_in(46,58) <= s_locks_lower_out(47,58);

		normal_cell_46_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,59),
			fetch              => s_fetch(46,59),
			data_in            => s_data_in(46,59),
			data_out           => s_data_out(46,59),
			out1               => s_out1(46,59),
			out2               => s_out2(46,59),
			lock_lower_row_out => s_locks_lower_out(46,59),
			lock_lower_row_in  => s_locks_lower_in(46,59),
			in1                => s_in1(46,59),
			in2                => s_in2(46,59),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(59)
		);
	s_in1(46,59)            <= s_out1(47,59);
	s_in2(46,59)            <= s_out2(47,60);
	s_locks_lower_in(46,59) <= s_locks_lower_out(47,59);

		last_col_cell_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(46,60),
			fetch              => s_fetch(46,60),
			data_in            => s_data_in(46,60),
			data_out           => s_data_out(46,60),
			out1               => s_out1(46,60),
			out2               => s_out2(46,60),
			lock_lower_row_out => s_locks_lower_out(46,60),
			lock_lower_row_in  => s_locks_lower_in(46,60),
			in1                => s_in1(46,60),
			in2                => (others => '0'),
			lock_row           => s_locks(46),
			piv_found          => s_piv_found,
			row_data           => s_row_data(46),
			col_data           => s_col_data(60)
		);
	s_in1(46,60)            <= s_out1(47,60);
	s_locks_lower_in(46,60) <= s_locks_lower_out(47,60);

		normal_cell_47_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,1),
			fetch              => s_fetch(47,1),
			data_in            => s_data_in(47,1),
			data_out           => s_data_out(47,1),
			out1               => s_out1(47,1),
			out2               => s_out2(47,1),
			lock_lower_row_out => s_locks_lower_out(47,1),
			lock_lower_row_in  => s_locks_lower_in(47,1),
			in1                => s_in1(47,1),
			in2                => s_in2(47,1),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(1)
		);
	s_in1(47,1)            <= s_out1(48,1);
	s_in2(47,1)            <= s_out2(48,2);
	s_locks_lower_in(47,1) <= s_locks_lower_out(48,1);

		normal_cell_47_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,2),
			fetch              => s_fetch(47,2),
			data_in            => s_data_in(47,2),
			data_out           => s_data_out(47,2),
			out1               => s_out1(47,2),
			out2               => s_out2(47,2),
			lock_lower_row_out => s_locks_lower_out(47,2),
			lock_lower_row_in  => s_locks_lower_in(47,2),
			in1                => s_in1(47,2),
			in2                => s_in2(47,2),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(2)
		);
	s_in1(47,2)            <= s_out1(48,2);
	s_in2(47,2)            <= s_out2(48,3);
	s_locks_lower_in(47,2) <= s_locks_lower_out(48,2);

		normal_cell_47_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,3),
			fetch              => s_fetch(47,3),
			data_in            => s_data_in(47,3),
			data_out           => s_data_out(47,3),
			out1               => s_out1(47,3),
			out2               => s_out2(47,3),
			lock_lower_row_out => s_locks_lower_out(47,3),
			lock_lower_row_in  => s_locks_lower_in(47,3),
			in1                => s_in1(47,3),
			in2                => s_in2(47,3),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(3)
		);
	s_in1(47,3)            <= s_out1(48,3);
	s_in2(47,3)            <= s_out2(48,4);
	s_locks_lower_in(47,3) <= s_locks_lower_out(48,3);

		normal_cell_47_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,4),
			fetch              => s_fetch(47,4),
			data_in            => s_data_in(47,4),
			data_out           => s_data_out(47,4),
			out1               => s_out1(47,4),
			out2               => s_out2(47,4),
			lock_lower_row_out => s_locks_lower_out(47,4),
			lock_lower_row_in  => s_locks_lower_in(47,4),
			in1                => s_in1(47,4),
			in2                => s_in2(47,4),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(4)
		);
	s_in1(47,4)            <= s_out1(48,4);
	s_in2(47,4)            <= s_out2(48,5);
	s_locks_lower_in(47,4) <= s_locks_lower_out(48,4);

		normal_cell_47_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,5),
			fetch              => s_fetch(47,5),
			data_in            => s_data_in(47,5),
			data_out           => s_data_out(47,5),
			out1               => s_out1(47,5),
			out2               => s_out2(47,5),
			lock_lower_row_out => s_locks_lower_out(47,5),
			lock_lower_row_in  => s_locks_lower_in(47,5),
			in1                => s_in1(47,5),
			in2                => s_in2(47,5),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(5)
		);
	s_in1(47,5)            <= s_out1(48,5);
	s_in2(47,5)            <= s_out2(48,6);
	s_locks_lower_in(47,5) <= s_locks_lower_out(48,5);

		normal_cell_47_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,6),
			fetch              => s_fetch(47,6),
			data_in            => s_data_in(47,6),
			data_out           => s_data_out(47,6),
			out1               => s_out1(47,6),
			out2               => s_out2(47,6),
			lock_lower_row_out => s_locks_lower_out(47,6),
			lock_lower_row_in  => s_locks_lower_in(47,6),
			in1                => s_in1(47,6),
			in2                => s_in2(47,6),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(6)
		);
	s_in1(47,6)            <= s_out1(48,6);
	s_in2(47,6)            <= s_out2(48,7);
	s_locks_lower_in(47,6) <= s_locks_lower_out(48,6);

		normal_cell_47_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,7),
			fetch              => s_fetch(47,7),
			data_in            => s_data_in(47,7),
			data_out           => s_data_out(47,7),
			out1               => s_out1(47,7),
			out2               => s_out2(47,7),
			lock_lower_row_out => s_locks_lower_out(47,7),
			lock_lower_row_in  => s_locks_lower_in(47,7),
			in1                => s_in1(47,7),
			in2                => s_in2(47,7),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(7)
		);
	s_in1(47,7)            <= s_out1(48,7);
	s_in2(47,7)            <= s_out2(48,8);
	s_locks_lower_in(47,7) <= s_locks_lower_out(48,7);

		normal_cell_47_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,8),
			fetch              => s_fetch(47,8),
			data_in            => s_data_in(47,8),
			data_out           => s_data_out(47,8),
			out1               => s_out1(47,8),
			out2               => s_out2(47,8),
			lock_lower_row_out => s_locks_lower_out(47,8),
			lock_lower_row_in  => s_locks_lower_in(47,8),
			in1                => s_in1(47,8),
			in2                => s_in2(47,8),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(8)
		);
	s_in1(47,8)            <= s_out1(48,8);
	s_in2(47,8)            <= s_out2(48,9);
	s_locks_lower_in(47,8) <= s_locks_lower_out(48,8);

		normal_cell_47_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,9),
			fetch              => s_fetch(47,9),
			data_in            => s_data_in(47,9),
			data_out           => s_data_out(47,9),
			out1               => s_out1(47,9),
			out2               => s_out2(47,9),
			lock_lower_row_out => s_locks_lower_out(47,9),
			lock_lower_row_in  => s_locks_lower_in(47,9),
			in1                => s_in1(47,9),
			in2                => s_in2(47,9),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(9)
		);
	s_in1(47,9)            <= s_out1(48,9);
	s_in2(47,9)            <= s_out2(48,10);
	s_locks_lower_in(47,9) <= s_locks_lower_out(48,9);

		normal_cell_47_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,10),
			fetch              => s_fetch(47,10),
			data_in            => s_data_in(47,10),
			data_out           => s_data_out(47,10),
			out1               => s_out1(47,10),
			out2               => s_out2(47,10),
			lock_lower_row_out => s_locks_lower_out(47,10),
			lock_lower_row_in  => s_locks_lower_in(47,10),
			in1                => s_in1(47,10),
			in2                => s_in2(47,10),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(10)
		);
	s_in1(47,10)            <= s_out1(48,10);
	s_in2(47,10)            <= s_out2(48,11);
	s_locks_lower_in(47,10) <= s_locks_lower_out(48,10);

		normal_cell_47_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,11),
			fetch              => s_fetch(47,11),
			data_in            => s_data_in(47,11),
			data_out           => s_data_out(47,11),
			out1               => s_out1(47,11),
			out2               => s_out2(47,11),
			lock_lower_row_out => s_locks_lower_out(47,11),
			lock_lower_row_in  => s_locks_lower_in(47,11),
			in1                => s_in1(47,11),
			in2                => s_in2(47,11),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(11)
		);
	s_in1(47,11)            <= s_out1(48,11);
	s_in2(47,11)            <= s_out2(48,12);
	s_locks_lower_in(47,11) <= s_locks_lower_out(48,11);

		normal_cell_47_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,12),
			fetch              => s_fetch(47,12),
			data_in            => s_data_in(47,12),
			data_out           => s_data_out(47,12),
			out1               => s_out1(47,12),
			out2               => s_out2(47,12),
			lock_lower_row_out => s_locks_lower_out(47,12),
			lock_lower_row_in  => s_locks_lower_in(47,12),
			in1                => s_in1(47,12),
			in2                => s_in2(47,12),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(12)
		);
	s_in1(47,12)            <= s_out1(48,12);
	s_in2(47,12)            <= s_out2(48,13);
	s_locks_lower_in(47,12) <= s_locks_lower_out(48,12);

		normal_cell_47_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,13),
			fetch              => s_fetch(47,13),
			data_in            => s_data_in(47,13),
			data_out           => s_data_out(47,13),
			out1               => s_out1(47,13),
			out2               => s_out2(47,13),
			lock_lower_row_out => s_locks_lower_out(47,13),
			lock_lower_row_in  => s_locks_lower_in(47,13),
			in1                => s_in1(47,13),
			in2                => s_in2(47,13),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(13)
		);
	s_in1(47,13)            <= s_out1(48,13);
	s_in2(47,13)            <= s_out2(48,14);
	s_locks_lower_in(47,13) <= s_locks_lower_out(48,13);

		normal_cell_47_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,14),
			fetch              => s_fetch(47,14),
			data_in            => s_data_in(47,14),
			data_out           => s_data_out(47,14),
			out1               => s_out1(47,14),
			out2               => s_out2(47,14),
			lock_lower_row_out => s_locks_lower_out(47,14),
			lock_lower_row_in  => s_locks_lower_in(47,14),
			in1                => s_in1(47,14),
			in2                => s_in2(47,14),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(14)
		);
	s_in1(47,14)            <= s_out1(48,14);
	s_in2(47,14)            <= s_out2(48,15);
	s_locks_lower_in(47,14) <= s_locks_lower_out(48,14);

		normal_cell_47_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,15),
			fetch              => s_fetch(47,15),
			data_in            => s_data_in(47,15),
			data_out           => s_data_out(47,15),
			out1               => s_out1(47,15),
			out2               => s_out2(47,15),
			lock_lower_row_out => s_locks_lower_out(47,15),
			lock_lower_row_in  => s_locks_lower_in(47,15),
			in1                => s_in1(47,15),
			in2                => s_in2(47,15),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(15)
		);
	s_in1(47,15)            <= s_out1(48,15);
	s_in2(47,15)            <= s_out2(48,16);
	s_locks_lower_in(47,15) <= s_locks_lower_out(48,15);

		normal_cell_47_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,16),
			fetch              => s_fetch(47,16),
			data_in            => s_data_in(47,16),
			data_out           => s_data_out(47,16),
			out1               => s_out1(47,16),
			out2               => s_out2(47,16),
			lock_lower_row_out => s_locks_lower_out(47,16),
			lock_lower_row_in  => s_locks_lower_in(47,16),
			in1                => s_in1(47,16),
			in2                => s_in2(47,16),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(16)
		);
	s_in1(47,16)            <= s_out1(48,16);
	s_in2(47,16)            <= s_out2(48,17);
	s_locks_lower_in(47,16) <= s_locks_lower_out(48,16);

		normal_cell_47_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,17),
			fetch              => s_fetch(47,17),
			data_in            => s_data_in(47,17),
			data_out           => s_data_out(47,17),
			out1               => s_out1(47,17),
			out2               => s_out2(47,17),
			lock_lower_row_out => s_locks_lower_out(47,17),
			lock_lower_row_in  => s_locks_lower_in(47,17),
			in1                => s_in1(47,17),
			in2                => s_in2(47,17),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(17)
		);
	s_in1(47,17)            <= s_out1(48,17);
	s_in2(47,17)            <= s_out2(48,18);
	s_locks_lower_in(47,17) <= s_locks_lower_out(48,17);

		normal_cell_47_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,18),
			fetch              => s_fetch(47,18),
			data_in            => s_data_in(47,18),
			data_out           => s_data_out(47,18),
			out1               => s_out1(47,18),
			out2               => s_out2(47,18),
			lock_lower_row_out => s_locks_lower_out(47,18),
			lock_lower_row_in  => s_locks_lower_in(47,18),
			in1                => s_in1(47,18),
			in2                => s_in2(47,18),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(18)
		);
	s_in1(47,18)            <= s_out1(48,18);
	s_in2(47,18)            <= s_out2(48,19);
	s_locks_lower_in(47,18) <= s_locks_lower_out(48,18);

		normal_cell_47_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,19),
			fetch              => s_fetch(47,19),
			data_in            => s_data_in(47,19),
			data_out           => s_data_out(47,19),
			out1               => s_out1(47,19),
			out2               => s_out2(47,19),
			lock_lower_row_out => s_locks_lower_out(47,19),
			lock_lower_row_in  => s_locks_lower_in(47,19),
			in1                => s_in1(47,19),
			in2                => s_in2(47,19),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(19)
		);
	s_in1(47,19)            <= s_out1(48,19);
	s_in2(47,19)            <= s_out2(48,20);
	s_locks_lower_in(47,19) <= s_locks_lower_out(48,19);

		normal_cell_47_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,20),
			fetch              => s_fetch(47,20),
			data_in            => s_data_in(47,20),
			data_out           => s_data_out(47,20),
			out1               => s_out1(47,20),
			out2               => s_out2(47,20),
			lock_lower_row_out => s_locks_lower_out(47,20),
			lock_lower_row_in  => s_locks_lower_in(47,20),
			in1                => s_in1(47,20),
			in2                => s_in2(47,20),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(20)
		);
	s_in1(47,20)            <= s_out1(48,20);
	s_in2(47,20)            <= s_out2(48,21);
	s_locks_lower_in(47,20) <= s_locks_lower_out(48,20);

		normal_cell_47_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,21),
			fetch              => s_fetch(47,21),
			data_in            => s_data_in(47,21),
			data_out           => s_data_out(47,21),
			out1               => s_out1(47,21),
			out2               => s_out2(47,21),
			lock_lower_row_out => s_locks_lower_out(47,21),
			lock_lower_row_in  => s_locks_lower_in(47,21),
			in1                => s_in1(47,21),
			in2                => s_in2(47,21),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(21)
		);
	s_in1(47,21)            <= s_out1(48,21);
	s_in2(47,21)            <= s_out2(48,22);
	s_locks_lower_in(47,21) <= s_locks_lower_out(48,21);

		normal_cell_47_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,22),
			fetch              => s_fetch(47,22),
			data_in            => s_data_in(47,22),
			data_out           => s_data_out(47,22),
			out1               => s_out1(47,22),
			out2               => s_out2(47,22),
			lock_lower_row_out => s_locks_lower_out(47,22),
			lock_lower_row_in  => s_locks_lower_in(47,22),
			in1                => s_in1(47,22),
			in2                => s_in2(47,22),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(22)
		);
	s_in1(47,22)            <= s_out1(48,22);
	s_in2(47,22)            <= s_out2(48,23);
	s_locks_lower_in(47,22) <= s_locks_lower_out(48,22);

		normal_cell_47_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,23),
			fetch              => s_fetch(47,23),
			data_in            => s_data_in(47,23),
			data_out           => s_data_out(47,23),
			out1               => s_out1(47,23),
			out2               => s_out2(47,23),
			lock_lower_row_out => s_locks_lower_out(47,23),
			lock_lower_row_in  => s_locks_lower_in(47,23),
			in1                => s_in1(47,23),
			in2                => s_in2(47,23),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(23)
		);
	s_in1(47,23)            <= s_out1(48,23);
	s_in2(47,23)            <= s_out2(48,24);
	s_locks_lower_in(47,23) <= s_locks_lower_out(48,23);

		normal_cell_47_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,24),
			fetch              => s_fetch(47,24),
			data_in            => s_data_in(47,24),
			data_out           => s_data_out(47,24),
			out1               => s_out1(47,24),
			out2               => s_out2(47,24),
			lock_lower_row_out => s_locks_lower_out(47,24),
			lock_lower_row_in  => s_locks_lower_in(47,24),
			in1                => s_in1(47,24),
			in2                => s_in2(47,24),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(24)
		);
	s_in1(47,24)            <= s_out1(48,24);
	s_in2(47,24)            <= s_out2(48,25);
	s_locks_lower_in(47,24) <= s_locks_lower_out(48,24);

		normal_cell_47_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,25),
			fetch              => s_fetch(47,25),
			data_in            => s_data_in(47,25),
			data_out           => s_data_out(47,25),
			out1               => s_out1(47,25),
			out2               => s_out2(47,25),
			lock_lower_row_out => s_locks_lower_out(47,25),
			lock_lower_row_in  => s_locks_lower_in(47,25),
			in1                => s_in1(47,25),
			in2                => s_in2(47,25),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(25)
		);
	s_in1(47,25)            <= s_out1(48,25);
	s_in2(47,25)            <= s_out2(48,26);
	s_locks_lower_in(47,25) <= s_locks_lower_out(48,25);

		normal_cell_47_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,26),
			fetch              => s_fetch(47,26),
			data_in            => s_data_in(47,26),
			data_out           => s_data_out(47,26),
			out1               => s_out1(47,26),
			out2               => s_out2(47,26),
			lock_lower_row_out => s_locks_lower_out(47,26),
			lock_lower_row_in  => s_locks_lower_in(47,26),
			in1                => s_in1(47,26),
			in2                => s_in2(47,26),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(26)
		);
	s_in1(47,26)            <= s_out1(48,26);
	s_in2(47,26)            <= s_out2(48,27);
	s_locks_lower_in(47,26) <= s_locks_lower_out(48,26);

		normal_cell_47_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,27),
			fetch              => s_fetch(47,27),
			data_in            => s_data_in(47,27),
			data_out           => s_data_out(47,27),
			out1               => s_out1(47,27),
			out2               => s_out2(47,27),
			lock_lower_row_out => s_locks_lower_out(47,27),
			lock_lower_row_in  => s_locks_lower_in(47,27),
			in1                => s_in1(47,27),
			in2                => s_in2(47,27),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(27)
		);
	s_in1(47,27)            <= s_out1(48,27);
	s_in2(47,27)            <= s_out2(48,28);
	s_locks_lower_in(47,27) <= s_locks_lower_out(48,27);

		normal_cell_47_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,28),
			fetch              => s_fetch(47,28),
			data_in            => s_data_in(47,28),
			data_out           => s_data_out(47,28),
			out1               => s_out1(47,28),
			out2               => s_out2(47,28),
			lock_lower_row_out => s_locks_lower_out(47,28),
			lock_lower_row_in  => s_locks_lower_in(47,28),
			in1                => s_in1(47,28),
			in2                => s_in2(47,28),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(28)
		);
	s_in1(47,28)            <= s_out1(48,28);
	s_in2(47,28)            <= s_out2(48,29);
	s_locks_lower_in(47,28) <= s_locks_lower_out(48,28);

		normal_cell_47_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,29),
			fetch              => s_fetch(47,29),
			data_in            => s_data_in(47,29),
			data_out           => s_data_out(47,29),
			out1               => s_out1(47,29),
			out2               => s_out2(47,29),
			lock_lower_row_out => s_locks_lower_out(47,29),
			lock_lower_row_in  => s_locks_lower_in(47,29),
			in1                => s_in1(47,29),
			in2                => s_in2(47,29),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(29)
		);
	s_in1(47,29)            <= s_out1(48,29);
	s_in2(47,29)            <= s_out2(48,30);
	s_locks_lower_in(47,29) <= s_locks_lower_out(48,29);

		normal_cell_47_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,30),
			fetch              => s_fetch(47,30),
			data_in            => s_data_in(47,30),
			data_out           => s_data_out(47,30),
			out1               => s_out1(47,30),
			out2               => s_out2(47,30),
			lock_lower_row_out => s_locks_lower_out(47,30),
			lock_lower_row_in  => s_locks_lower_in(47,30),
			in1                => s_in1(47,30),
			in2                => s_in2(47,30),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(30)
		);
	s_in1(47,30)            <= s_out1(48,30);
	s_in2(47,30)            <= s_out2(48,31);
	s_locks_lower_in(47,30) <= s_locks_lower_out(48,30);

		normal_cell_47_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,31),
			fetch              => s_fetch(47,31),
			data_in            => s_data_in(47,31),
			data_out           => s_data_out(47,31),
			out1               => s_out1(47,31),
			out2               => s_out2(47,31),
			lock_lower_row_out => s_locks_lower_out(47,31),
			lock_lower_row_in  => s_locks_lower_in(47,31),
			in1                => s_in1(47,31),
			in2                => s_in2(47,31),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(31)
		);
	s_in1(47,31)            <= s_out1(48,31);
	s_in2(47,31)            <= s_out2(48,32);
	s_locks_lower_in(47,31) <= s_locks_lower_out(48,31);

		normal_cell_47_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,32),
			fetch              => s_fetch(47,32),
			data_in            => s_data_in(47,32),
			data_out           => s_data_out(47,32),
			out1               => s_out1(47,32),
			out2               => s_out2(47,32),
			lock_lower_row_out => s_locks_lower_out(47,32),
			lock_lower_row_in  => s_locks_lower_in(47,32),
			in1                => s_in1(47,32),
			in2                => s_in2(47,32),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(32)
		);
	s_in1(47,32)            <= s_out1(48,32);
	s_in2(47,32)            <= s_out2(48,33);
	s_locks_lower_in(47,32) <= s_locks_lower_out(48,32);

		normal_cell_47_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,33),
			fetch              => s_fetch(47,33),
			data_in            => s_data_in(47,33),
			data_out           => s_data_out(47,33),
			out1               => s_out1(47,33),
			out2               => s_out2(47,33),
			lock_lower_row_out => s_locks_lower_out(47,33),
			lock_lower_row_in  => s_locks_lower_in(47,33),
			in1                => s_in1(47,33),
			in2                => s_in2(47,33),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(33)
		);
	s_in1(47,33)            <= s_out1(48,33);
	s_in2(47,33)            <= s_out2(48,34);
	s_locks_lower_in(47,33) <= s_locks_lower_out(48,33);

		normal_cell_47_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,34),
			fetch              => s_fetch(47,34),
			data_in            => s_data_in(47,34),
			data_out           => s_data_out(47,34),
			out1               => s_out1(47,34),
			out2               => s_out2(47,34),
			lock_lower_row_out => s_locks_lower_out(47,34),
			lock_lower_row_in  => s_locks_lower_in(47,34),
			in1                => s_in1(47,34),
			in2                => s_in2(47,34),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(34)
		);
	s_in1(47,34)            <= s_out1(48,34);
	s_in2(47,34)            <= s_out2(48,35);
	s_locks_lower_in(47,34) <= s_locks_lower_out(48,34);

		normal_cell_47_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,35),
			fetch              => s_fetch(47,35),
			data_in            => s_data_in(47,35),
			data_out           => s_data_out(47,35),
			out1               => s_out1(47,35),
			out2               => s_out2(47,35),
			lock_lower_row_out => s_locks_lower_out(47,35),
			lock_lower_row_in  => s_locks_lower_in(47,35),
			in1                => s_in1(47,35),
			in2                => s_in2(47,35),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(35)
		);
	s_in1(47,35)            <= s_out1(48,35);
	s_in2(47,35)            <= s_out2(48,36);
	s_locks_lower_in(47,35) <= s_locks_lower_out(48,35);

		normal_cell_47_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,36),
			fetch              => s_fetch(47,36),
			data_in            => s_data_in(47,36),
			data_out           => s_data_out(47,36),
			out1               => s_out1(47,36),
			out2               => s_out2(47,36),
			lock_lower_row_out => s_locks_lower_out(47,36),
			lock_lower_row_in  => s_locks_lower_in(47,36),
			in1                => s_in1(47,36),
			in2                => s_in2(47,36),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(36)
		);
	s_in1(47,36)            <= s_out1(48,36);
	s_in2(47,36)            <= s_out2(48,37);
	s_locks_lower_in(47,36) <= s_locks_lower_out(48,36);

		normal_cell_47_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,37),
			fetch              => s_fetch(47,37),
			data_in            => s_data_in(47,37),
			data_out           => s_data_out(47,37),
			out1               => s_out1(47,37),
			out2               => s_out2(47,37),
			lock_lower_row_out => s_locks_lower_out(47,37),
			lock_lower_row_in  => s_locks_lower_in(47,37),
			in1                => s_in1(47,37),
			in2                => s_in2(47,37),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(37)
		);
	s_in1(47,37)            <= s_out1(48,37);
	s_in2(47,37)            <= s_out2(48,38);
	s_locks_lower_in(47,37) <= s_locks_lower_out(48,37);

		normal_cell_47_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,38),
			fetch              => s_fetch(47,38),
			data_in            => s_data_in(47,38),
			data_out           => s_data_out(47,38),
			out1               => s_out1(47,38),
			out2               => s_out2(47,38),
			lock_lower_row_out => s_locks_lower_out(47,38),
			lock_lower_row_in  => s_locks_lower_in(47,38),
			in1                => s_in1(47,38),
			in2                => s_in2(47,38),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(38)
		);
	s_in1(47,38)            <= s_out1(48,38);
	s_in2(47,38)            <= s_out2(48,39);
	s_locks_lower_in(47,38) <= s_locks_lower_out(48,38);

		normal_cell_47_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,39),
			fetch              => s_fetch(47,39),
			data_in            => s_data_in(47,39),
			data_out           => s_data_out(47,39),
			out1               => s_out1(47,39),
			out2               => s_out2(47,39),
			lock_lower_row_out => s_locks_lower_out(47,39),
			lock_lower_row_in  => s_locks_lower_in(47,39),
			in1                => s_in1(47,39),
			in2                => s_in2(47,39),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(39)
		);
	s_in1(47,39)            <= s_out1(48,39);
	s_in2(47,39)            <= s_out2(48,40);
	s_locks_lower_in(47,39) <= s_locks_lower_out(48,39);

		normal_cell_47_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,40),
			fetch              => s_fetch(47,40),
			data_in            => s_data_in(47,40),
			data_out           => s_data_out(47,40),
			out1               => s_out1(47,40),
			out2               => s_out2(47,40),
			lock_lower_row_out => s_locks_lower_out(47,40),
			lock_lower_row_in  => s_locks_lower_in(47,40),
			in1                => s_in1(47,40),
			in2                => s_in2(47,40),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(40)
		);
	s_in1(47,40)            <= s_out1(48,40);
	s_in2(47,40)            <= s_out2(48,41);
	s_locks_lower_in(47,40) <= s_locks_lower_out(48,40);

		normal_cell_47_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,41),
			fetch              => s_fetch(47,41),
			data_in            => s_data_in(47,41),
			data_out           => s_data_out(47,41),
			out1               => s_out1(47,41),
			out2               => s_out2(47,41),
			lock_lower_row_out => s_locks_lower_out(47,41),
			lock_lower_row_in  => s_locks_lower_in(47,41),
			in1                => s_in1(47,41),
			in2                => s_in2(47,41),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(41)
		);
	s_in1(47,41)            <= s_out1(48,41);
	s_in2(47,41)            <= s_out2(48,42);
	s_locks_lower_in(47,41) <= s_locks_lower_out(48,41);

		normal_cell_47_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,42),
			fetch              => s_fetch(47,42),
			data_in            => s_data_in(47,42),
			data_out           => s_data_out(47,42),
			out1               => s_out1(47,42),
			out2               => s_out2(47,42),
			lock_lower_row_out => s_locks_lower_out(47,42),
			lock_lower_row_in  => s_locks_lower_in(47,42),
			in1                => s_in1(47,42),
			in2                => s_in2(47,42),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(42)
		);
	s_in1(47,42)            <= s_out1(48,42);
	s_in2(47,42)            <= s_out2(48,43);
	s_locks_lower_in(47,42) <= s_locks_lower_out(48,42);

		normal_cell_47_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,43),
			fetch              => s_fetch(47,43),
			data_in            => s_data_in(47,43),
			data_out           => s_data_out(47,43),
			out1               => s_out1(47,43),
			out2               => s_out2(47,43),
			lock_lower_row_out => s_locks_lower_out(47,43),
			lock_lower_row_in  => s_locks_lower_in(47,43),
			in1                => s_in1(47,43),
			in2                => s_in2(47,43),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(43)
		);
	s_in1(47,43)            <= s_out1(48,43);
	s_in2(47,43)            <= s_out2(48,44);
	s_locks_lower_in(47,43) <= s_locks_lower_out(48,43);

		normal_cell_47_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,44),
			fetch              => s_fetch(47,44),
			data_in            => s_data_in(47,44),
			data_out           => s_data_out(47,44),
			out1               => s_out1(47,44),
			out2               => s_out2(47,44),
			lock_lower_row_out => s_locks_lower_out(47,44),
			lock_lower_row_in  => s_locks_lower_in(47,44),
			in1                => s_in1(47,44),
			in2                => s_in2(47,44),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(44)
		);
	s_in1(47,44)            <= s_out1(48,44);
	s_in2(47,44)            <= s_out2(48,45);
	s_locks_lower_in(47,44) <= s_locks_lower_out(48,44);

		normal_cell_47_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,45),
			fetch              => s_fetch(47,45),
			data_in            => s_data_in(47,45),
			data_out           => s_data_out(47,45),
			out1               => s_out1(47,45),
			out2               => s_out2(47,45),
			lock_lower_row_out => s_locks_lower_out(47,45),
			lock_lower_row_in  => s_locks_lower_in(47,45),
			in1                => s_in1(47,45),
			in2                => s_in2(47,45),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(45)
		);
	s_in1(47,45)            <= s_out1(48,45);
	s_in2(47,45)            <= s_out2(48,46);
	s_locks_lower_in(47,45) <= s_locks_lower_out(48,45);

		normal_cell_47_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,46),
			fetch              => s_fetch(47,46),
			data_in            => s_data_in(47,46),
			data_out           => s_data_out(47,46),
			out1               => s_out1(47,46),
			out2               => s_out2(47,46),
			lock_lower_row_out => s_locks_lower_out(47,46),
			lock_lower_row_in  => s_locks_lower_in(47,46),
			in1                => s_in1(47,46),
			in2                => s_in2(47,46),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(46)
		);
	s_in1(47,46)            <= s_out1(48,46);
	s_in2(47,46)            <= s_out2(48,47);
	s_locks_lower_in(47,46) <= s_locks_lower_out(48,46);

		normal_cell_47_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,47),
			fetch              => s_fetch(47,47),
			data_in            => s_data_in(47,47),
			data_out           => s_data_out(47,47),
			out1               => s_out1(47,47),
			out2               => s_out2(47,47),
			lock_lower_row_out => s_locks_lower_out(47,47),
			lock_lower_row_in  => s_locks_lower_in(47,47),
			in1                => s_in1(47,47),
			in2                => s_in2(47,47),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(47)
		);
	s_in1(47,47)            <= s_out1(48,47);
	s_in2(47,47)            <= s_out2(48,48);
	s_locks_lower_in(47,47) <= s_locks_lower_out(48,47);

		normal_cell_47_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,48),
			fetch              => s_fetch(47,48),
			data_in            => s_data_in(47,48),
			data_out           => s_data_out(47,48),
			out1               => s_out1(47,48),
			out2               => s_out2(47,48),
			lock_lower_row_out => s_locks_lower_out(47,48),
			lock_lower_row_in  => s_locks_lower_in(47,48),
			in1                => s_in1(47,48),
			in2                => s_in2(47,48),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(48)
		);
	s_in1(47,48)            <= s_out1(48,48);
	s_in2(47,48)            <= s_out2(48,49);
	s_locks_lower_in(47,48) <= s_locks_lower_out(48,48);

		normal_cell_47_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,49),
			fetch              => s_fetch(47,49),
			data_in            => s_data_in(47,49),
			data_out           => s_data_out(47,49),
			out1               => s_out1(47,49),
			out2               => s_out2(47,49),
			lock_lower_row_out => s_locks_lower_out(47,49),
			lock_lower_row_in  => s_locks_lower_in(47,49),
			in1                => s_in1(47,49),
			in2                => s_in2(47,49),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(49)
		);
	s_in1(47,49)            <= s_out1(48,49);
	s_in2(47,49)            <= s_out2(48,50);
	s_locks_lower_in(47,49) <= s_locks_lower_out(48,49);

		normal_cell_47_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,50),
			fetch              => s_fetch(47,50),
			data_in            => s_data_in(47,50),
			data_out           => s_data_out(47,50),
			out1               => s_out1(47,50),
			out2               => s_out2(47,50),
			lock_lower_row_out => s_locks_lower_out(47,50),
			lock_lower_row_in  => s_locks_lower_in(47,50),
			in1                => s_in1(47,50),
			in2                => s_in2(47,50),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(50)
		);
	s_in1(47,50)            <= s_out1(48,50);
	s_in2(47,50)            <= s_out2(48,51);
	s_locks_lower_in(47,50) <= s_locks_lower_out(48,50);

		normal_cell_47_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,51),
			fetch              => s_fetch(47,51),
			data_in            => s_data_in(47,51),
			data_out           => s_data_out(47,51),
			out1               => s_out1(47,51),
			out2               => s_out2(47,51),
			lock_lower_row_out => s_locks_lower_out(47,51),
			lock_lower_row_in  => s_locks_lower_in(47,51),
			in1                => s_in1(47,51),
			in2                => s_in2(47,51),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(51)
		);
	s_in1(47,51)            <= s_out1(48,51);
	s_in2(47,51)            <= s_out2(48,52);
	s_locks_lower_in(47,51) <= s_locks_lower_out(48,51);

		normal_cell_47_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,52),
			fetch              => s_fetch(47,52),
			data_in            => s_data_in(47,52),
			data_out           => s_data_out(47,52),
			out1               => s_out1(47,52),
			out2               => s_out2(47,52),
			lock_lower_row_out => s_locks_lower_out(47,52),
			lock_lower_row_in  => s_locks_lower_in(47,52),
			in1                => s_in1(47,52),
			in2                => s_in2(47,52),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(52)
		);
	s_in1(47,52)            <= s_out1(48,52);
	s_in2(47,52)            <= s_out2(48,53);
	s_locks_lower_in(47,52) <= s_locks_lower_out(48,52);

		normal_cell_47_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,53),
			fetch              => s_fetch(47,53),
			data_in            => s_data_in(47,53),
			data_out           => s_data_out(47,53),
			out1               => s_out1(47,53),
			out2               => s_out2(47,53),
			lock_lower_row_out => s_locks_lower_out(47,53),
			lock_lower_row_in  => s_locks_lower_in(47,53),
			in1                => s_in1(47,53),
			in2                => s_in2(47,53),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(53)
		);
	s_in1(47,53)            <= s_out1(48,53);
	s_in2(47,53)            <= s_out2(48,54);
	s_locks_lower_in(47,53) <= s_locks_lower_out(48,53);

		normal_cell_47_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,54),
			fetch              => s_fetch(47,54),
			data_in            => s_data_in(47,54),
			data_out           => s_data_out(47,54),
			out1               => s_out1(47,54),
			out2               => s_out2(47,54),
			lock_lower_row_out => s_locks_lower_out(47,54),
			lock_lower_row_in  => s_locks_lower_in(47,54),
			in1                => s_in1(47,54),
			in2                => s_in2(47,54),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(54)
		);
	s_in1(47,54)            <= s_out1(48,54);
	s_in2(47,54)            <= s_out2(48,55);
	s_locks_lower_in(47,54) <= s_locks_lower_out(48,54);

		normal_cell_47_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,55),
			fetch              => s_fetch(47,55),
			data_in            => s_data_in(47,55),
			data_out           => s_data_out(47,55),
			out1               => s_out1(47,55),
			out2               => s_out2(47,55),
			lock_lower_row_out => s_locks_lower_out(47,55),
			lock_lower_row_in  => s_locks_lower_in(47,55),
			in1                => s_in1(47,55),
			in2                => s_in2(47,55),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(55)
		);
	s_in1(47,55)            <= s_out1(48,55);
	s_in2(47,55)            <= s_out2(48,56);
	s_locks_lower_in(47,55) <= s_locks_lower_out(48,55);

		normal_cell_47_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,56),
			fetch              => s_fetch(47,56),
			data_in            => s_data_in(47,56),
			data_out           => s_data_out(47,56),
			out1               => s_out1(47,56),
			out2               => s_out2(47,56),
			lock_lower_row_out => s_locks_lower_out(47,56),
			lock_lower_row_in  => s_locks_lower_in(47,56),
			in1                => s_in1(47,56),
			in2                => s_in2(47,56),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(56)
		);
	s_in1(47,56)            <= s_out1(48,56);
	s_in2(47,56)            <= s_out2(48,57);
	s_locks_lower_in(47,56) <= s_locks_lower_out(48,56);

		normal_cell_47_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,57),
			fetch              => s_fetch(47,57),
			data_in            => s_data_in(47,57),
			data_out           => s_data_out(47,57),
			out1               => s_out1(47,57),
			out2               => s_out2(47,57),
			lock_lower_row_out => s_locks_lower_out(47,57),
			lock_lower_row_in  => s_locks_lower_in(47,57),
			in1                => s_in1(47,57),
			in2                => s_in2(47,57),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(57)
		);
	s_in1(47,57)            <= s_out1(48,57);
	s_in2(47,57)            <= s_out2(48,58);
	s_locks_lower_in(47,57) <= s_locks_lower_out(48,57);

		normal_cell_47_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,58),
			fetch              => s_fetch(47,58),
			data_in            => s_data_in(47,58),
			data_out           => s_data_out(47,58),
			out1               => s_out1(47,58),
			out2               => s_out2(47,58),
			lock_lower_row_out => s_locks_lower_out(47,58),
			lock_lower_row_in  => s_locks_lower_in(47,58),
			in1                => s_in1(47,58),
			in2                => s_in2(47,58),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(58)
		);
	s_in1(47,58)            <= s_out1(48,58);
	s_in2(47,58)            <= s_out2(48,59);
	s_locks_lower_in(47,58) <= s_locks_lower_out(48,58);

		normal_cell_47_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,59),
			fetch              => s_fetch(47,59),
			data_in            => s_data_in(47,59),
			data_out           => s_data_out(47,59),
			out1               => s_out1(47,59),
			out2               => s_out2(47,59),
			lock_lower_row_out => s_locks_lower_out(47,59),
			lock_lower_row_in  => s_locks_lower_in(47,59),
			in1                => s_in1(47,59),
			in2                => s_in2(47,59),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(59)
		);
	s_in1(47,59)            <= s_out1(48,59);
	s_in2(47,59)            <= s_out2(48,60);
	s_locks_lower_in(47,59) <= s_locks_lower_out(48,59);

		last_col_cell_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(47,60),
			fetch              => s_fetch(47,60),
			data_in            => s_data_in(47,60),
			data_out           => s_data_out(47,60),
			out1               => s_out1(47,60),
			out2               => s_out2(47,60),
			lock_lower_row_out => s_locks_lower_out(47,60),
			lock_lower_row_in  => s_locks_lower_in(47,60),
			in1                => s_in1(47,60),
			in2                => (others => '0'),
			lock_row           => s_locks(47),
			piv_found          => s_piv_found,
			row_data           => s_row_data(47),
			col_data           => s_col_data(60)
		);
	s_in1(47,60)            <= s_out1(48,60);
	s_locks_lower_in(47,60) <= s_locks_lower_out(48,60);

		normal_cell_48_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,1),
			fetch              => s_fetch(48,1),
			data_in            => s_data_in(48,1),
			data_out           => s_data_out(48,1),
			out1               => s_out1(48,1),
			out2               => s_out2(48,1),
			lock_lower_row_out => s_locks_lower_out(48,1),
			lock_lower_row_in  => s_locks_lower_in(48,1),
			in1                => s_in1(48,1),
			in2                => s_in2(48,1),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(1)
		);
	s_in1(48,1)            <= s_out1(49,1);
	s_in2(48,1)            <= s_out2(49,2);
	s_locks_lower_in(48,1) <= s_locks_lower_out(49,1);

		normal_cell_48_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,2),
			fetch              => s_fetch(48,2),
			data_in            => s_data_in(48,2),
			data_out           => s_data_out(48,2),
			out1               => s_out1(48,2),
			out2               => s_out2(48,2),
			lock_lower_row_out => s_locks_lower_out(48,2),
			lock_lower_row_in  => s_locks_lower_in(48,2),
			in1                => s_in1(48,2),
			in2                => s_in2(48,2),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(2)
		);
	s_in1(48,2)            <= s_out1(49,2);
	s_in2(48,2)            <= s_out2(49,3);
	s_locks_lower_in(48,2) <= s_locks_lower_out(49,2);

		normal_cell_48_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,3),
			fetch              => s_fetch(48,3),
			data_in            => s_data_in(48,3),
			data_out           => s_data_out(48,3),
			out1               => s_out1(48,3),
			out2               => s_out2(48,3),
			lock_lower_row_out => s_locks_lower_out(48,3),
			lock_lower_row_in  => s_locks_lower_in(48,3),
			in1                => s_in1(48,3),
			in2                => s_in2(48,3),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(3)
		);
	s_in1(48,3)            <= s_out1(49,3);
	s_in2(48,3)            <= s_out2(49,4);
	s_locks_lower_in(48,3) <= s_locks_lower_out(49,3);

		normal_cell_48_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,4),
			fetch              => s_fetch(48,4),
			data_in            => s_data_in(48,4),
			data_out           => s_data_out(48,4),
			out1               => s_out1(48,4),
			out2               => s_out2(48,4),
			lock_lower_row_out => s_locks_lower_out(48,4),
			lock_lower_row_in  => s_locks_lower_in(48,4),
			in1                => s_in1(48,4),
			in2                => s_in2(48,4),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(4)
		);
	s_in1(48,4)            <= s_out1(49,4);
	s_in2(48,4)            <= s_out2(49,5);
	s_locks_lower_in(48,4) <= s_locks_lower_out(49,4);

		normal_cell_48_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,5),
			fetch              => s_fetch(48,5),
			data_in            => s_data_in(48,5),
			data_out           => s_data_out(48,5),
			out1               => s_out1(48,5),
			out2               => s_out2(48,5),
			lock_lower_row_out => s_locks_lower_out(48,5),
			lock_lower_row_in  => s_locks_lower_in(48,5),
			in1                => s_in1(48,5),
			in2                => s_in2(48,5),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(5)
		);
	s_in1(48,5)            <= s_out1(49,5);
	s_in2(48,5)            <= s_out2(49,6);
	s_locks_lower_in(48,5) <= s_locks_lower_out(49,5);

		normal_cell_48_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,6),
			fetch              => s_fetch(48,6),
			data_in            => s_data_in(48,6),
			data_out           => s_data_out(48,6),
			out1               => s_out1(48,6),
			out2               => s_out2(48,6),
			lock_lower_row_out => s_locks_lower_out(48,6),
			lock_lower_row_in  => s_locks_lower_in(48,6),
			in1                => s_in1(48,6),
			in2                => s_in2(48,6),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(6)
		);
	s_in1(48,6)            <= s_out1(49,6);
	s_in2(48,6)            <= s_out2(49,7);
	s_locks_lower_in(48,6) <= s_locks_lower_out(49,6);

		normal_cell_48_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,7),
			fetch              => s_fetch(48,7),
			data_in            => s_data_in(48,7),
			data_out           => s_data_out(48,7),
			out1               => s_out1(48,7),
			out2               => s_out2(48,7),
			lock_lower_row_out => s_locks_lower_out(48,7),
			lock_lower_row_in  => s_locks_lower_in(48,7),
			in1                => s_in1(48,7),
			in2                => s_in2(48,7),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(7)
		);
	s_in1(48,7)            <= s_out1(49,7);
	s_in2(48,7)            <= s_out2(49,8);
	s_locks_lower_in(48,7) <= s_locks_lower_out(49,7);

		normal_cell_48_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,8),
			fetch              => s_fetch(48,8),
			data_in            => s_data_in(48,8),
			data_out           => s_data_out(48,8),
			out1               => s_out1(48,8),
			out2               => s_out2(48,8),
			lock_lower_row_out => s_locks_lower_out(48,8),
			lock_lower_row_in  => s_locks_lower_in(48,8),
			in1                => s_in1(48,8),
			in2                => s_in2(48,8),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(8)
		);
	s_in1(48,8)            <= s_out1(49,8);
	s_in2(48,8)            <= s_out2(49,9);
	s_locks_lower_in(48,8) <= s_locks_lower_out(49,8);

		normal_cell_48_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,9),
			fetch              => s_fetch(48,9),
			data_in            => s_data_in(48,9),
			data_out           => s_data_out(48,9),
			out1               => s_out1(48,9),
			out2               => s_out2(48,9),
			lock_lower_row_out => s_locks_lower_out(48,9),
			lock_lower_row_in  => s_locks_lower_in(48,9),
			in1                => s_in1(48,9),
			in2                => s_in2(48,9),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(9)
		);
	s_in1(48,9)            <= s_out1(49,9);
	s_in2(48,9)            <= s_out2(49,10);
	s_locks_lower_in(48,9) <= s_locks_lower_out(49,9);

		normal_cell_48_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,10),
			fetch              => s_fetch(48,10),
			data_in            => s_data_in(48,10),
			data_out           => s_data_out(48,10),
			out1               => s_out1(48,10),
			out2               => s_out2(48,10),
			lock_lower_row_out => s_locks_lower_out(48,10),
			lock_lower_row_in  => s_locks_lower_in(48,10),
			in1                => s_in1(48,10),
			in2                => s_in2(48,10),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(10)
		);
	s_in1(48,10)            <= s_out1(49,10);
	s_in2(48,10)            <= s_out2(49,11);
	s_locks_lower_in(48,10) <= s_locks_lower_out(49,10);

		normal_cell_48_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,11),
			fetch              => s_fetch(48,11),
			data_in            => s_data_in(48,11),
			data_out           => s_data_out(48,11),
			out1               => s_out1(48,11),
			out2               => s_out2(48,11),
			lock_lower_row_out => s_locks_lower_out(48,11),
			lock_lower_row_in  => s_locks_lower_in(48,11),
			in1                => s_in1(48,11),
			in2                => s_in2(48,11),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(11)
		);
	s_in1(48,11)            <= s_out1(49,11);
	s_in2(48,11)            <= s_out2(49,12);
	s_locks_lower_in(48,11) <= s_locks_lower_out(49,11);

		normal_cell_48_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,12),
			fetch              => s_fetch(48,12),
			data_in            => s_data_in(48,12),
			data_out           => s_data_out(48,12),
			out1               => s_out1(48,12),
			out2               => s_out2(48,12),
			lock_lower_row_out => s_locks_lower_out(48,12),
			lock_lower_row_in  => s_locks_lower_in(48,12),
			in1                => s_in1(48,12),
			in2                => s_in2(48,12),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(12)
		);
	s_in1(48,12)            <= s_out1(49,12);
	s_in2(48,12)            <= s_out2(49,13);
	s_locks_lower_in(48,12) <= s_locks_lower_out(49,12);

		normal_cell_48_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,13),
			fetch              => s_fetch(48,13),
			data_in            => s_data_in(48,13),
			data_out           => s_data_out(48,13),
			out1               => s_out1(48,13),
			out2               => s_out2(48,13),
			lock_lower_row_out => s_locks_lower_out(48,13),
			lock_lower_row_in  => s_locks_lower_in(48,13),
			in1                => s_in1(48,13),
			in2                => s_in2(48,13),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(13)
		);
	s_in1(48,13)            <= s_out1(49,13);
	s_in2(48,13)            <= s_out2(49,14);
	s_locks_lower_in(48,13) <= s_locks_lower_out(49,13);

		normal_cell_48_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,14),
			fetch              => s_fetch(48,14),
			data_in            => s_data_in(48,14),
			data_out           => s_data_out(48,14),
			out1               => s_out1(48,14),
			out2               => s_out2(48,14),
			lock_lower_row_out => s_locks_lower_out(48,14),
			lock_lower_row_in  => s_locks_lower_in(48,14),
			in1                => s_in1(48,14),
			in2                => s_in2(48,14),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(14)
		);
	s_in1(48,14)            <= s_out1(49,14);
	s_in2(48,14)            <= s_out2(49,15);
	s_locks_lower_in(48,14) <= s_locks_lower_out(49,14);

		normal_cell_48_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,15),
			fetch              => s_fetch(48,15),
			data_in            => s_data_in(48,15),
			data_out           => s_data_out(48,15),
			out1               => s_out1(48,15),
			out2               => s_out2(48,15),
			lock_lower_row_out => s_locks_lower_out(48,15),
			lock_lower_row_in  => s_locks_lower_in(48,15),
			in1                => s_in1(48,15),
			in2                => s_in2(48,15),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(15)
		);
	s_in1(48,15)            <= s_out1(49,15);
	s_in2(48,15)            <= s_out2(49,16);
	s_locks_lower_in(48,15) <= s_locks_lower_out(49,15);

		normal_cell_48_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,16),
			fetch              => s_fetch(48,16),
			data_in            => s_data_in(48,16),
			data_out           => s_data_out(48,16),
			out1               => s_out1(48,16),
			out2               => s_out2(48,16),
			lock_lower_row_out => s_locks_lower_out(48,16),
			lock_lower_row_in  => s_locks_lower_in(48,16),
			in1                => s_in1(48,16),
			in2                => s_in2(48,16),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(16)
		);
	s_in1(48,16)            <= s_out1(49,16);
	s_in2(48,16)            <= s_out2(49,17);
	s_locks_lower_in(48,16) <= s_locks_lower_out(49,16);

		normal_cell_48_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,17),
			fetch              => s_fetch(48,17),
			data_in            => s_data_in(48,17),
			data_out           => s_data_out(48,17),
			out1               => s_out1(48,17),
			out2               => s_out2(48,17),
			lock_lower_row_out => s_locks_lower_out(48,17),
			lock_lower_row_in  => s_locks_lower_in(48,17),
			in1                => s_in1(48,17),
			in2                => s_in2(48,17),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(17)
		);
	s_in1(48,17)            <= s_out1(49,17);
	s_in2(48,17)            <= s_out2(49,18);
	s_locks_lower_in(48,17) <= s_locks_lower_out(49,17);

		normal_cell_48_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,18),
			fetch              => s_fetch(48,18),
			data_in            => s_data_in(48,18),
			data_out           => s_data_out(48,18),
			out1               => s_out1(48,18),
			out2               => s_out2(48,18),
			lock_lower_row_out => s_locks_lower_out(48,18),
			lock_lower_row_in  => s_locks_lower_in(48,18),
			in1                => s_in1(48,18),
			in2                => s_in2(48,18),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(18)
		);
	s_in1(48,18)            <= s_out1(49,18);
	s_in2(48,18)            <= s_out2(49,19);
	s_locks_lower_in(48,18) <= s_locks_lower_out(49,18);

		normal_cell_48_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,19),
			fetch              => s_fetch(48,19),
			data_in            => s_data_in(48,19),
			data_out           => s_data_out(48,19),
			out1               => s_out1(48,19),
			out2               => s_out2(48,19),
			lock_lower_row_out => s_locks_lower_out(48,19),
			lock_lower_row_in  => s_locks_lower_in(48,19),
			in1                => s_in1(48,19),
			in2                => s_in2(48,19),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(19)
		);
	s_in1(48,19)            <= s_out1(49,19);
	s_in2(48,19)            <= s_out2(49,20);
	s_locks_lower_in(48,19) <= s_locks_lower_out(49,19);

		normal_cell_48_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,20),
			fetch              => s_fetch(48,20),
			data_in            => s_data_in(48,20),
			data_out           => s_data_out(48,20),
			out1               => s_out1(48,20),
			out2               => s_out2(48,20),
			lock_lower_row_out => s_locks_lower_out(48,20),
			lock_lower_row_in  => s_locks_lower_in(48,20),
			in1                => s_in1(48,20),
			in2                => s_in2(48,20),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(20)
		);
	s_in1(48,20)            <= s_out1(49,20);
	s_in2(48,20)            <= s_out2(49,21);
	s_locks_lower_in(48,20) <= s_locks_lower_out(49,20);

		normal_cell_48_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,21),
			fetch              => s_fetch(48,21),
			data_in            => s_data_in(48,21),
			data_out           => s_data_out(48,21),
			out1               => s_out1(48,21),
			out2               => s_out2(48,21),
			lock_lower_row_out => s_locks_lower_out(48,21),
			lock_lower_row_in  => s_locks_lower_in(48,21),
			in1                => s_in1(48,21),
			in2                => s_in2(48,21),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(21)
		);
	s_in1(48,21)            <= s_out1(49,21);
	s_in2(48,21)            <= s_out2(49,22);
	s_locks_lower_in(48,21) <= s_locks_lower_out(49,21);

		normal_cell_48_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,22),
			fetch              => s_fetch(48,22),
			data_in            => s_data_in(48,22),
			data_out           => s_data_out(48,22),
			out1               => s_out1(48,22),
			out2               => s_out2(48,22),
			lock_lower_row_out => s_locks_lower_out(48,22),
			lock_lower_row_in  => s_locks_lower_in(48,22),
			in1                => s_in1(48,22),
			in2                => s_in2(48,22),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(22)
		);
	s_in1(48,22)            <= s_out1(49,22);
	s_in2(48,22)            <= s_out2(49,23);
	s_locks_lower_in(48,22) <= s_locks_lower_out(49,22);

		normal_cell_48_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,23),
			fetch              => s_fetch(48,23),
			data_in            => s_data_in(48,23),
			data_out           => s_data_out(48,23),
			out1               => s_out1(48,23),
			out2               => s_out2(48,23),
			lock_lower_row_out => s_locks_lower_out(48,23),
			lock_lower_row_in  => s_locks_lower_in(48,23),
			in1                => s_in1(48,23),
			in2                => s_in2(48,23),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(23)
		);
	s_in1(48,23)            <= s_out1(49,23);
	s_in2(48,23)            <= s_out2(49,24);
	s_locks_lower_in(48,23) <= s_locks_lower_out(49,23);

		normal_cell_48_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,24),
			fetch              => s_fetch(48,24),
			data_in            => s_data_in(48,24),
			data_out           => s_data_out(48,24),
			out1               => s_out1(48,24),
			out2               => s_out2(48,24),
			lock_lower_row_out => s_locks_lower_out(48,24),
			lock_lower_row_in  => s_locks_lower_in(48,24),
			in1                => s_in1(48,24),
			in2                => s_in2(48,24),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(24)
		);
	s_in1(48,24)            <= s_out1(49,24);
	s_in2(48,24)            <= s_out2(49,25);
	s_locks_lower_in(48,24) <= s_locks_lower_out(49,24);

		normal_cell_48_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,25),
			fetch              => s_fetch(48,25),
			data_in            => s_data_in(48,25),
			data_out           => s_data_out(48,25),
			out1               => s_out1(48,25),
			out2               => s_out2(48,25),
			lock_lower_row_out => s_locks_lower_out(48,25),
			lock_lower_row_in  => s_locks_lower_in(48,25),
			in1                => s_in1(48,25),
			in2                => s_in2(48,25),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(25)
		);
	s_in1(48,25)            <= s_out1(49,25);
	s_in2(48,25)            <= s_out2(49,26);
	s_locks_lower_in(48,25) <= s_locks_lower_out(49,25);

		normal_cell_48_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,26),
			fetch              => s_fetch(48,26),
			data_in            => s_data_in(48,26),
			data_out           => s_data_out(48,26),
			out1               => s_out1(48,26),
			out2               => s_out2(48,26),
			lock_lower_row_out => s_locks_lower_out(48,26),
			lock_lower_row_in  => s_locks_lower_in(48,26),
			in1                => s_in1(48,26),
			in2                => s_in2(48,26),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(26)
		);
	s_in1(48,26)            <= s_out1(49,26);
	s_in2(48,26)            <= s_out2(49,27);
	s_locks_lower_in(48,26) <= s_locks_lower_out(49,26);

		normal_cell_48_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,27),
			fetch              => s_fetch(48,27),
			data_in            => s_data_in(48,27),
			data_out           => s_data_out(48,27),
			out1               => s_out1(48,27),
			out2               => s_out2(48,27),
			lock_lower_row_out => s_locks_lower_out(48,27),
			lock_lower_row_in  => s_locks_lower_in(48,27),
			in1                => s_in1(48,27),
			in2                => s_in2(48,27),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(27)
		);
	s_in1(48,27)            <= s_out1(49,27);
	s_in2(48,27)            <= s_out2(49,28);
	s_locks_lower_in(48,27) <= s_locks_lower_out(49,27);

		normal_cell_48_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,28),
			fetch              => s_fetch(48,28),
			data_in            => s_data_in(48,28),
			data_out           => s_data_out(48,28),
			out1               => s_out1(48,28),
			out2               => s_out2(48,28),
			lock_lower_row_out => s_locks_lower_out(48,28),
			lock_lower_row_in  => s_locks_lower_in(48,28),
			in1                => s_in1(48,28),
			in2                => s_in2(48,28),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(28)
		);
	s_in1(48,28)            <= s_out1(49,28);
	s_in2(48,28)            <= s_out2(49,29);
	s_locks_lower_in(48,28) <= s_locks_lower_out(49,28);

		normal_cell_48_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,29),
			fetch              => s_fetch(48,29),
			data_in            => s_data_in(48,29),
			data_out           => s_data_out(48,29),
			out1               => s_out1(48,29),
			out2               => s_out2(48,29),
			lock_lower_row_out => s_locks_lower_out(48,29),
			lock_lower_row_in  => s_locks_lower_in(48,29),
			in1                => s_in1(48,29),
			in2                => s_in2(48,29),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(29)
		);
	s_in1(48,29)            <= s_out1(49,29);
	s_in2(48,29)            <= s_out2(49,30);
	s_locks_lower_in(48,29) <= s_locks_lower_out(49,29);

		normal_cell_48_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,30),
			fetch              => s_fetch(48,30),
			data_in            => s_data_in(48,30),
			data_out           => s_data_out(48,30),
			out1               => s_out1(48,30),
			out2               => s_out2(48,30),
			lock_lower_row_out => s_locks_lower_out(48,30),
			lock_lower_row_in  => s_locks_lower_in(48,30),
			in1                => s_in1(48,30),
			in2                => s_in2(48,30),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(30)
		);
	s_in1(48,30)            <= s_out1(49,30);
	s_in2(48,30)            <= s_out2(49,31);
	s_locks_lower_in(48,30) <= s_locks_lower_out(49,30);

		normal_cell_48_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,31),
			fetch              => s_fetch(48,31),
			data_in            => s_data_in(48,31),
			data_out           => s_data_out(48,31),
			out1               => s_out1(48,31),
			out2               => s_out2(48,31),
			lock_lower_row_out => s_locks_lower_out(48,31),
			lock_lower_row_in  => s_locks_lower_in(48,31),
			in1                => s_in1(48,31),
			in2                => s_in2(48,31),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(31)
		);
	s_in1(48,31)            <= s_out1(49,31);
	s_in2(48,31)            <= s_out2(49,32);
	s_locks_lower_in(48,31) <= s_locks_lower_out(49,31);

		normal_cell_48_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,32),
			fetch              => s_fetch(48,32),
			data_in            => s_data_in(48,32),
			data_out           => s_data_out(48,32),
			out1               => s_out1(48,32),
			out2               => s_out2(48,32),
			lock_lower_row_out => s_locks_lower_out(48,32),
			lock_lower_row_in  => s_locks_lower_in(48,32),
			in1                => s_in1(48,32),
			in2                => s_in2(48,32),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(32)
		);
	s_in1(48,32)            <= s_out1(49,32);
	s_in2(48,32)            <= s_out2(49,33);
	s_locks_lower_in(48,32) <= s_locks_lower_out(49,32);

		normal_cell_48_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,33),
			fetch              => s_fetch(48,33),
			data_in            => s_data_in(48,33),
			data_out           => s_data_out(48,33),
			out1               => s_out1(48,33),
			out2               => s_out2(48,33),
			lock_lower_row_out => s_locks_lower_out(48,33),
			lock_lower_row_in  => s_locks_lower_in(48,33),
			in1                => s_in1(48,33),
			in2                => s_in2(48,33),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(33)
		);
	s_in1(48,33)            <= s_out1(49,33);
	s_in2(48,33)            <= s_out2(49,34);
	s_locks_lower_in(48,33) <= s_locks_lower_out(49,33);

		normal_cell_48_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,34),
			fetch              => s_fetch(48,34),
			data_in            => s_data_in(48,34),
			data_out           => s_data_out(48,34),
			out1               => s_out1(48,34),
			out2               => s_out2(48,34),
			lock_lower_row_out => s_locks_lower_out(48,34),
			lock_lower_row_in  => s_locks_lower_in(48,34),
			in1                => s_in1(48,34),
			in2                => s_in2(48,34),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(34)
		);
	s_in1(48,34)            <= s_out1(49,34);
	s_in2(48,34)            <= s_out2(49,35);
	s_locks_lower_in(48,34) <= s_locks_lower_out(49,34);

		normal_cell_48_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,35),
			fetch              => s_fetch(48,35),
			data_in            => s_data_in(48,35),
			data_out           => s_data_out(48,35),
			out1               => s_out1(48,35),
			out2               => s_out2(48,35),
			lock_lower_row_out => s_locks_lower_out(48,35),
			lock_lower_row_in  => s_locks_lower_in(48,35),
			in1                => s_in1(48,35),
			in2                => s_in2(48,35),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(35)
		);
	s_in1(48,35)            <= s_out1(49,35);
	s_in2(48,35)            <= s_out2(49,36);
	s_locks_lower_in(48,35) <= s_locks_lower_out(49,35);

		normal_cell_48_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,36),
			fetch              => s_fetch(48,36),
			data_in            => s_data_in(48,36),
			data_out           => s_data_out(48,36),
			out1               => s_out1(48,36),
			out2               => s_out2(48,36),
			lock_lower_row_out => s_locks_lower_out(48,36),
			lock_lower_row_in  => s_locks_lower_in(48,36),
			in1                => s_in1(48,36),
			in2                => s_in2(48,36),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(36)
		);
	s_in1(48,36)            <= s_out1(49,36);
	s_in2(48,36)            <= s_out2(49,37);
	s_locks_lower_in(48,36) <= s_locks_lower_out(49,36);

		normal_cell_48_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,37),
			fetch              => s_fetch(48,37),
			data_in            => s_data_in(48,37),
			data_out           => s_data_out(48,37),
			out1               => s_out1(48,37),
			out2               => s_out2(48,37),
			lock_lower_row_out => s_locks_lower_out(48,37),
			lock_lower_row_in  => s_locks_lower_in(48,37),
			in1                => s_in1(48,37),
			in2                => s_in2(48,37),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(37)
		);
	s_in1(48,37)            <= s_out1(49,37);
	s_in2(48,37)            <= s_out2(49,38);
	s_locks_lower_in(48,37) <= s_locks_lower_out(49,37);

		normal_cell_48_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,38),
			fetch              => s_fetch(48,38),
			data_in            => s_data_in(48,38),
			data_out           => s_data_out(48,38),
			out1               => s_out1(48,38),
			out2               => s_out2(48,38),
			lock_lower_row_out => s_locks_lower_out(48,38),
			lock_lower_row_in  => s_locks_lower_in(48,38),
			in1                => s_in1(48,38),
			in2                => s_in2(48,38),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(38)
		);
	s_in1(48,38)            <= s_out1(49,38);
	s_in2(48,38)            <= s_out2(49,39);
	s_locks_lower_in(48,38) <= s_locks_lower_out(49,38);

		normal_cell_48_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,39),
			fetch              => s_fetch(48,39),
			data_in            => s_data_in(48,39),
			data_out           => s_data_out(48,39),
			out1               => s_out1(48,39),
			out2               => s_out2(48,39),
			lock_lower_row_out => s_locks_lower_out(48,39),
			lock_lower_row_in  => s_locks_lower_in(48,39),
			in1                => s_in1(48,39),
			in2                => s_in2(48,39),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(39)
		);
	s_in1(48,39)            <= s_out1(49,39);
	s_in2(48,39)            <= s_out2(49,40);
	s_locks_lower_in(48,39) <= s_locks_lower_out(49,39);

		normal_cell_48_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,40),
			fetch              => s_fetch(48,40),
			data_in            => s_data_in(48,40),
			data_out           => s_data_out(48,40),
			out1               => s_out1(48,40),
			out2               => s_out2(48,40),
			lock_lower_row_out => s_locks_lower_out(48,40),
			lock_lower_row_in  => s_locks_lower_in(48,40),
			in1                => s_in1(48,40),
			in2                => s_in2(48,40),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(40)
		);
	s_in1(48,40)            <= s_out1(49,40);
	s_in2(48,40)            <= s_out2(49,41);
	s_locks_lower_in(48,40) <= s_locks_lower_out(49,40);

		normal_cell_48_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,41),
			fetch              => s_fetch(48,41),
			data_in            => s_data_in(48,41),
			data_out           => s_data_out(48,41),
			out1               => s_out1(48,41),
			out2               => s_out2(48,41),
			lock_lower_row_out => s_locks_lower_out(48,41),
			lock_lower_row_in  => s_locks_lower_in(48,41),
			in1                => s_in1(48,41),
			in2                => s_in2(48,41),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(41)
		);
	s_in1(48,41)            <= s_out1(49,41);
	s_in2(48,41)            <= s_out2(49,42);
	s_locks_lower_in(48,41) <= s_locks_lower_out(49,41);

		normal_cell_48_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,42),
			fetch              => s_fetch(48,42),
			data_in            => s_data_in(48,42),
			data_out           => s_data_out(48,42),
			out1               => s_out1(48,42),
			out2               => s_out2(48,42),
			lock_lower_row_out => s_locks_lower_out(48,42),
			lock_lower_row_in  => s_locks_lower_in(48,42),
			in1                => s_in1(48,42),
			in2                => s_in2(48,42),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(42)
		);
	s_in1(48,42)            <= s_out1(49,42);
	s_in2(48,42)            <= s_out2(49,43);
	s_locks_lower_in(48,42) <= s_locks_lower_out(49,42);

		normal_cell_48_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,43),
			fetch              => s_fetch(48,43),
			data_in            => s_data_in(48,43),
			data_out           => s_data_out(48,43),
			out1               => s_out1(48,43),
			out2               => s_out2(48,43),
			lock_lower_row_out => s_locks_lower_out(48,43),
			lock_lower_row_in  => s_locks_lower_in(48,43),
			in1                => s_in1(48,43),
			in2                => s_in2(48,43),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(43)
		);
	s_in1(48,43)            <= s_out1(49,43);
	s_in2(48,43)            <= s_out2(49,44);
	s_locks_lower_in(48,43) <= s_locks_lower_out(49,43);

		normal_cell_48_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,44),
			fetch              => s_fetch(48,44),
			data_in            => s_data_in(48,44),
			data_out           => s_data_out(48,44),
			out1               => s_out1(48,44),
			out2               => s_out2(48,44),
			lock_lower_row_out => s_locks_lower_out(48,44),
			lock_lower_row_in  => s_locks_lower_in(48,44),
			in1                => s_in1(48,44),
			in2                => s_in2(48,44),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(44)
		);
	s_in1(48,44)            <= s_out1(49,44);
	s_in2(48,44)            <= s_out2(49,45);
	s_locks_lower_in(48,44) <= s_locks_lower_out(49,44);

		normal_cell_48_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,45),
			fetch              => s_fetch(48,45),
			data_in            => s_data_in(48,45),
			data_out           => s_data_out(48,45),
			out1               => s_out1(48,45),
			out2               => s_out2(48,45),
			lock_lower_row_out => s_locks_lower_out(48,45),
			lock_lower_row_in  => s_locks_lower_in(48,45),
			in1                => s_in1(48,45),
			in2                => s_in2(48,45),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(45)
		);
	s_in1(48,45)            <= s_out1(49,45);
	s_in2(48,45)            <= s_out2(49,46);
	s_locks_lower_in(48,45) <= s_locks_lower_out(49,45);

		normal_cell_48_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,46),
			fetch              => s_fetch(48,46),
			data_in            => s_data_in(48,46),
			data_out           => s_data_out(48,46),
			out1               => s_out1(48,46),
			out2               => s_out2(48,46),
			lock_lower_row_out => s_locks_lower_out(48,46),
			lock_lower_row_in  => s_locks_lower_in(48,46),
			in1                => s_in1(48,46),
			in2                => s_in2(48,46),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(46)
		);
	s_in1(48,46)            <= s_out1(49,46);
	s_in2(48,46)            <= s_out2(49,47);
	s_locks_lower_in(48,46) <= s_locks_lower_out(49,46);

		normal_cell_48_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,47),
			fetch              => s_fetch(48,47),
			data_in            => s_data_in(48,47),
			data_out           => s_data_out(48,47),
			out1               => s_out1(48,47),
			out2               => s_out2(48,47),
			lock_lower_row_out => s_locks_lower_out(48,47),
			lock_lower_row_in  => s_locks_lower_in(48,47),
			in1                => s_in1(48,47),
			in2                => s_in2(48,47),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(47)
		);
	s_in1(48,47)            <= s_out1(49,47);
	s_in2(48,47)            <= s_out2(49,48);
	s_locks_lower_in(48,47) <= s_locks_lower_out(49,47);

		normal_cell_48_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,48),
			fetch              => s_fetch(48,48),
			data_in            => s_data_in(48,48),
			data_out           => s_data_out(48,48),
			out1               => s_out1(48,48),
			out2               => s_out2(48,48),
			lock_lower_row_out => s_locks_lower_out(48,48),
			lock_lower_row_in  => s_locks_lower_in(48,48),
			in1                => s_in1(48,48),
			in2                => s_in2(48,48),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(48)
		);
	s_in1(48,48)            <= s_out1(49,48);
	s_in2(48,48)            <= s_out2(49,49);
	s_locks_lower_in(48,48) <= s_locks_lower_out(49,48);

		normal_cell_48_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,49),
			fetch              => s_fetch(48,49),
			data_in            => s_data_in(48,49),
			data_out           => s_data_out(48,49),
			out1               => s_out1(48,49),
			out2               => s_out2(48,49),
			lock_lower_row_out => s_locks_lower_out(48,49),
			lock_lower_row_in  => s_locks_lower_in(48,49),
			in1                => s_in1(48,49),
			in2                => s_in2(48,49),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(49)
		);
	s_in1(48,49)            <= s_out1(49,49);
	s_in2(48,49)            <= s_out2(49,50);
	s_locks_lower_in(48,49) <= s_locks_lower_out(49,49);

		normal_cell_48_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,50),
			fetch              => s_fetch(48,50),
			data_in            => s_data_in(48,50),
			data_out           => s_data_out(48,50),
			out1               => s_out1(48,50),
			out2               => s_out2(48,50),
			lock_lower_row_out => s_locks_lower_out(48,50),
			lock_lower_row_in  => s_locks_lower_in(48,50),
			in1                => s_in1(48,50),
			in2                => s_in2(48,50),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(50)
		);
	s_in1(48,50)            <= s_out1(49,50);
	s_in2(48,50)            <= s_out2(49,51);
	s_locks_lower_in(48,50) <= s_locks_lower_out(49,50);

		normal_cell_48_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,51),
			fetch              => s_fetch(48,51),
			data_in            => s_data_in(48,51),
			data_out           => s_data_out(48,51),
			out1               => s_out1(48,51),
			out2               => s_out2(48,51),
			lock_lower_row_out => s_locks_lower_out(48,51),
			lock_lower_row_in  => s_locks_lower_in(48,51),
			in1                => s_in1(48,51),
			in2                => s_in2(48,51),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(51)
		);
	s_in1(48,51)            <= s_out1(49,51);
	s_in2(48,51)            <= s_out2(49,52);
	s_locks_lower_in(48,51) <= s_locks_lower_out(49,51);

		normal_cell_48_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,52),
			fetch              => s_fetch(48,52),
			data_in            => s_data_in(48,52),
			data_out           => s_data_out(48,52),
			out1               => s_out1(48,52),
			out2               => s_out2(48,52),
			lock_lower_row_out => s_locks_lower_out(48,52),
			lock_lower_row_in  => s_locks_lower_in(48,52),
			in1                => s_in1(48,52),
			in2                => s_in2(48,52),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(52)
		);
	s_in1(48,52)            <= s_out1(49,52);
	s_in2(48,52)            <= s_out2(49,53);
	s_locks_lower_in(48,52) <= s_locks_lower_out(49,52);

		normal_cell_48_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,53),
			fetch              => s_fetch(48,53),
			data_in            => s_data_in(48,53),
			data_out           => s_data_out(48,53),
			out1               => s_out1(48,53),
			out2               => s_out2(48,53),
			lock_lower_row_out => s_locks_lower_out(48,53),
			lock_lower_row_in  => s_locks_lower_in(48,53),
			in1                => s_in1(48,53),
			in2                => s_in2(48,53),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(53)
		);
	s_in1(48,53)            <= s_out1(49,53);
	s_in2(48,53)            <= s_out2(49,54);
	s_locks_lower_in(48,53) <= s_locks_lower_out(49,53);

		normal_cell_48_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,54),
			fetch              => s_fetch(48,54),
			data_in            => s_data_in(48,54),
			data_out           => s_data_out(48,54),
			out1               => s_out1(48,54),
			out2               => s_out2(48,54),
			lock_lower_row_out => s_locks_lower_out(48,54),
			lock_lower_row_in  => s_locks_lower_in(48,54),
			in1                => s_in1(48,54),
			in2                => s_in2(48,54),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(54)
		);
	s_in1(48,54)            <= s_out1(49,54);
	s_in2(48,54)            <= s_out2(49,55);
	s_locks_lower_in(48,54) <= s_locks_lower_out(49,54);

		normal_cell_48_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,55),
			fetch              => s_fetch(48,55),
			data_in            => s_data_in(48,55),
			data_out           => s_data_out(48,55),
			out1               => s_out1(48,55),
			out2               => s_out2(48,55),
			lock_lower_row_out => s_locks_lower_out(48,55),
			lock_lower_row_in  => s_locks_lower_in(48,55),
			in1                => s_in1(48,55),
			in2                => s_in2(48,55),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(55)
		);
	s_in1(48,55)            <= s_out1(49,55);
	s_in2(48,55)            <= s_out2(49,56);
	s_locks_lower_in(48,55) <= s_locks_lower_out(49,55);

		normal_cell_48_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,56),
			fetch              => s_fetch(48,56),
			data_in            => s_data_in(48,56),
			data_out           => s_data_out(48,56),
			out1               => s_out1(48,56),
			out2               => s_out2(48,56),
			lock_lower_row_out => s_locks_lower_out(48,56),
			lock_lower_row_in  => s_locks_lower_in(48,56),
			in1                => s_in1(48,56),
			in2                => s_in2(48,56),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(56)
		);
	s_in1(48,56)            <= s_out1(49,56);
	s_in2(48,56)            <= s_out2(49,57);
	s_locks_lower_in(48,56) <= s_locks_lower_out(49,56);

		normal_cell_48_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,57),
			fetch              => s_fetch(48,57),
			data_in            => s_data_in(48,57),
			data_out           => s_data_out(48,57),
			out1               => s_out1(48,57),
			out2               => s_out2(48,57),
			lock_lower_row_out => s_locks_lower_out(48,57),
			lock_lower_row_in  => s_locks_lower_in(48,57),
			in1                => s_in1(48,57),
			in2                => s_in2(48,57),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(57)
		);
	s_in1(48,57)            <= s_out1(49,57);
	s_in2(48,57)            <= s_out2(49,58);
	s_locks_lower_in(48,57) <= s_locks_lower_out(49,57);

		normal_cell_48_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,58),
			fetch              => s_fetch(48,58),
			data_in            => s_data_in(48,58),
			data_out           => s_data_out(48,58),
			out1               => s_out1(48,58),
			out2               => s_out2(48,58),
			lock_lower_row_out => s_locks_lower_out(48,58),
			lock_lower_row_in  => s_locks_lower_in(48,58),
			in1                => s_in1(48,58),
			in2                => s_in2(48,58),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(58)
		);
	s_in1(48,58)            <= s_out1(49,58);
	s_in2(48,58)            <= s_out2(49,59);
	s_locks_lower_in(48,58) <= s_locks_lower_out(49,58);

		normal_cell_48_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,59),
			fetch              => s_fetch(48,59),
			data_in            => s_data_in(48,59),
			data_out           => s_data_out(48,59),
			out1               => s_out1(48,59),
			out2               => s_out2(48,59),
			lock_lower_row_out => s_locks_lower_out(48,59),
			lock_lower_row_in  => s_locks_lower_in(48,59),
			in1                => s_in1(48,59),
			in2                => s_in2(48,59),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(59)
		);
	s_in1(48,59)            <= s_out1(49,59);
	s_in2(48,59)            <= s_out2(49,60);
	s_locks_lower_in(48,59) <= s_locks_lower_out(49,59);

		last_col_cell_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(48,60),
			fetch              => s_fetch(48,60),
			data_in            => s_data_in(48,60),
			data_out           => s_data_out(48,60),
			out1               => s_out1(48,60),
			out2               => s_out2(48,60),
			lock_lower_row_out => s_locks_lower_out(48,60),
			lock_lower_row_in  => s_locks_lower_in(48,60),
			in1                => s_in1(48,60),
			in2                => (others => '0'),
			lock_row           => s_locks(48),
			piv_found          => s_piv_found,
			row_data           => s_row_data(48),
			col_data           => s_col_data(60)
		);
	s_in1(48,60)            <= s_out1(49,60);
	s_locks_lower_in(48,60) <= s_locks_lower_out(49,60);

		normal_cell_49_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,1),
			fetch              => s_fetch(49,1),
			data_in            => s_data_in(49,1),
			data_out           => s_data_out(49,1),
			out1               => s_out1(49,1),
			out2               => s_out2(49,1),
			lock_lower_row_out => s_locks_lower_out(49,1),
			lock_lower_row_in  => s_locks_lower_in(49,1),
			in1                => s_in1(49,1),
			in2                => s_in2(49,1),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(1)
		);
	s_in1(49,1)            <= s_out1(50,1);
	s_in2(49,1)            <= s_out2(50,2);
	s_locks_lower_in(49,1) <= s_locks_lower_out(50,1);

		normal_cell_49_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,2),
			fetch              => s_fetch(49,2),
			data_in            => s_data_in(49,2),
			data_out           => s_data_out(49,2),
			out1               => s_out1(49,2),
			out2               => s_out2(49,2),
			lock_lower_row_out => s_locks_lower_out(49,2),
			lock_lower_row_in  => s_locks_lower_in(49,2),
			in1                => s_in1(49,2),
			in2                => s_in2(49,2),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(2)
		);
	s_in1(49,2)            <= s_out1(50,2);
	s_in2(49,2)            <= s_out2(50,3);
	s_locks_lower_in(49,2) <= s_locks_lower_out(50,2);

		normal_cell_49_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,3),
			fetch              => s_fetch(49,3),
			data_in            => s_data_in(49,3),
			data_out           => s_data_out(49,3),
			out1               => s_out1(49,3),
			out2               => s_out2(49,3),
			lock_lower_row_out => s_locks_lower_out(49,3),
			lock_lower_row_in  => s_locks_lower_in(49,3),
			in1                => s_in1(49,3),
			in2                => s_in2(49,3),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(3)
		);
	s_in1(49,3)            <= s_out1(50,3);
	s_in2(49,3)            <= s_out2(50,4);
	s_locks_lower_in(49,3) <= s_locks_lower_out(50,3);

		normal_cell_49_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,4),
			fetch              => s_fetch(49,4),
			data_in            => s_data_in(49,4),
			data_out           => s_data_out(49,4),
			out1               => s_out1(49,4),
			out2               => s_out2(49,4),
			lock_lower_row_out => s_locks_lower_out(49,4),
			lock_lower_row_in  => s_locks_lower_in(49,4),
			in1                => s_in1(49,4),
			in2                => s_in2(49,4),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(4)
		);
	s_in1(49,4)            <= s_out1(50,4);
	s_in2(49,4)            <= s_out2(50,5);
	s_locks_lower_in(49,4) <= s_locks_lower_out(50,4);

		normal_cell_49_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,5),
			fetch              => s_fetch(49,5),
			data_in            => s_data_in(49,5),
			data_out           => s_data_out(49,5),
			out1               => s_out1(49,5),
			out2               => s_out2(49,5),
			lock_lower_row_out => s_locks_lower_out(49,5),
			lock_lower_row_in  => s_locks_lower_in(49,5),
			in1                => s_in1(49,5),
			in2                => s_in2(49,5),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(5)
		);
	s_in1(49,5)            <= s_out1(50,5);
	s_in2(49,5)            <= s_out2(50,6);
	s_locks_lower_in(49,5) <= s_locks_lower_out(50,5);

		normal_cell_49_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,6),
			fetch              => s_fetch(49,6),
			data_in            => s_data_in(49,6),
			data_out           => s_data_out(49,6),
			out1               => s_out1(49,6),
			out2               => s_out2(49,6),
			lock_lower_row_out => s_locks_lower_out(49,6),
			lock_lower_row_in  => s_locks_lower_in(49,6),
			in1                => s_in1(49,6),
			in2                => s_in2(49,6),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(6)
		);
	s_in1(49,6)            <= s_out1(50,6);
	s_in2(49,6)            <= s_out2(50,7);
	s_locks_lower_in(49,6) <= s_locks_lower_out(50,6);

		normal_cell_49_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,7),
			fetch              => s_fetch(49,7),
			data_in            => s_data_in(49,7),
			data_out           => s_data_out(49,7),
			out1               => s_out1(49,7),
			out2               => s_out2(49,7),
			lock_lower_row_out => s_locks_lower_out(49,7),
			lock_lower_row_in  => s_locks_lower_in(49,7),
			in1                => s_in1(49,7),
			in2                => s_in2(49,7),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(7)
		);
	s_in1(49,7)            <= s_out1(50,7);
	s_in2(49,7)            <= s_out2(50,8);
	s_locks_lower_in(49,7) <= s_locks_lower_out(50,7);

		normal_cell_49_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,8),
			fetch              => s_fetch(49,8),
			data_in            => s_data_in(49,8),
			data_out           => s_data_out(49,8),
			out1               => s_out1(49,8),
			out2               => s_out2(49,8),
			lock_lower_row_out => s_locks_lower_out(49,8),
			lock_lower_row_in  => s_locks_lower_in(49,8),
			in1                => s_in1(49,8),
			in2                => s_in2(49,8),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(8)
		);
	s_in1(49,8)            <= s_out1(50,8);
	s_in2(49,8)            <= s_out2(50,9);
	s_locks_lower_in(49,8) <= s_locks_lower_out(50,8);

		normal_cell_49_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,9),
			fetch              => s_fetch(49,9),
			data_in            => s_data_in(49,9),
			data_out           => s_data_out(49,9),
			out1               => s_out1(49,9),
			out2               => s_out2(49,9),
			lock_lower_row_out => s_locks_lower_out(49,9),
			lock_lower_row_in  => s_locks_lower_in(49,9),
			in1                => s_in1(49,9),
			in2                => s_in2(49,9),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(9)
		);
	s_in1(49,9)            <= s_out1(50,9);
	s_in2(49,9)            <= s_out2(50,10);
	s_locks_lower_in(49,9) <= s_locks_lower_out(50,9);

		normal_cell_49_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,10),
			fetch              => s_fetch(49,10),
			data_in            => s_data_in(49,10),
			data_out           => s_data_out(49,10),
			out1               => s_out1(49,10),
			out2               => s_out2(49,10),
			lock_lower_row_out => s_locks_lower_out(49,10),
			lock_lower_row_in  => s_locks_lower_in(49,10),
			in1                => s_in1(49,10),
			in2                => s_in2(49,10),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(10)
		);
	s_in1(49,10)            <= s_out1(50,10);
	s_in2(49,10)            <= s_out2(50,11);
	s_locks_lower_in(49,10) <= s_locks_lower_out(50,10);

		normal_cell_49_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,11),
			fetch              => s_fetch(49,11),
			data_in            => s_data_in(49,11),
			data_out           => s_data_out(49,11),
			out1               => s_out1(49,11),
			out2               => s_out2(49,11),
			lock_lower_row_out => s_locks_lower_out(49,11),
			lock_lower_row_in  => s_locks_lower_in(49,11),
			in1                => s_in1(49,11),
			in2                => s_in2(49,11),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(11)
		);
	s_in1(49,11)            <= s_out1(50,11);
	s_in2(49,11)            <= s_out2(50,12);
	s_locks_lower_in(49,11) <= s_locks_lower_out(50,11);

		normal_cell_49_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,12),
			fetch              => s_fetch(49,12),
			data_in            => s_data_in(49,12),
			data_out           => s_data_out(49,12),
			out1               => s_out1(49,12),
			out2               => s_out2(49,12),
			lock_lower_row_out => s_locks_lower_out(49,12),
			lock_lower_row_in  => s_locks_lower_in(49,12),
			in1                => s_in1(49,12),
			in2                => s_in2(49,12),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(12)
		);
	s_in1(49,12)            <= s_out1(50,12);
	s_in2(49,12)            <= s_out2(50,13);
	s_locks_lower_in(49,12) <= s_locks_lower_out(50,12);

		normal_cell_49_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,13),
			fetch              => s_fetch(49,13),
			data_in            => s_data_in(49,13),
			data_out           => s_data_out(49,13),
			out1               => s_out1(49,13),
			out2               => s_out2(49,13),
			lock_lower_row_out => s_locks_lower_out(49,13),
			lock_lower_row_in  => s_locks_lower_in(49,13),
			in1                => s_in1(49,13),
			in2                => s_in2(49,13),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(13)
		);
	s_in1(49,13)            <= s_out1(50,13);
	s_in2(49,13)            <= s_out2(50,14);
	s_locks_lower_in(49,13) <= s_locks_lower_out(50,13);

		normal_cell_49_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,14),
			fetch              => s_fetch(49,14),
			data_in            => s_data_in(49,14),
			data_out           => s_data_out(49,14),
			out1               => s_out1(49,14),
			out2               => s_out2(49,14),
			lock_lower_row_out => s_locks_lower_out(49,14),
			lock_lower_row_in  => s_locks_lower_in(49,14),
			in1                => s_in1(49,14),
			in2                => s_in2(49,14),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(14)
		);
	s_in1(49,14)            <= s_out1(50,14);
	s_in2(49,14)            <= s_out2(50,15);
	s_locks_lower_in(49,14) <= s_locks_lower_out(50,14);

		normal_cell_49_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,15),
			fetch              => s_fetch(49,15),
			data_in            => s_data_in(49,15),
			data_out           => s_data_out(49,15),
			out1               => s_out1(49,15),
			out2               => s_out2(49,15),
			lock_lower_row_out => s_locks_lower_out(49,15),
			lock_lower_row_in  => s_locks_lower_in(49,15),
			in1                => s_in1(49,15),
			in2                => s_in2(49,15),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(15)
		);
	s_in1(49,15)            <= s_out1(50,15);
	s_in2(49,15)            <= s_out2(50,16);
	s_locks_lower_in(49,15) <= s_locks_lower_out(50,15);

		normal_cell_49_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,16),
			fetch              => s_fetch(49,16),
			data_in            => s_data_in(49,16),
			data_out           => s_data_out(49,16),
			out1               => s_out1(49,16),
			out2               => s_out2(49,16),
			lock_lower_row_out => s_locks_lower_out(49,16),
			lock_lower_row_in  => s_locks_lower_in(49,16),
			in1                => s_in1(49,16),
			in2                => s_in2(49,16),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(16)
		);
	s_in1(49,16)            <= s_out1(50,16);
	s_in2(49,16)            <= s_out2(50,17);
	s_locks_lower_in(49,16) <= s_locks_lower_out(50,16);

		normal_cell_49_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,17),
			fetch              => s_fetch(49,17),
			data_in            => s_data_in(49,17),
			data_out           => s_data_out(49,17),
			out1               => s_out1(49,17),
			out2               => s_out2(49,17),
			lock_lower_row_out => s_locks_lower_out(49,17),
			lock_lower_row_in  => s_locks_lower_in(49,17),
			in1                => s_in1(49,17),
			in2                => s_in2(49,17),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(17)
		);
	s_in1(49,17)            <= s_out1(50,17);
	s_in2(49,17)            <= s_out2(50,18);
	s_locks_lower_in(49,17) <= s_locks_lower_out(50,17);

		normal_cell_49_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,18),
			fetch              => s_fetch(49,18),
			data_in            => s_data_in(49,18),
			data_out           => s_data_out(49,18),
			out1               => s_out1(49,18),
			out2               => s_out2(49,18),
			lock_lower_row_out => s_locks_lower_out(49,18),
			lock_lower_row_in  => s_locks_lower_in(49,18),
			in1                => s_in1(49,18),
			in2                => s_in2(49,18),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(18)
		);
	s_in1(49,18)            <= s_out1(50,18);
	s_in2(49,18)            <= s_out2(50,19);
	s_locks_lower_in(49,18) <= s_locks_lower_out(50,18);

		normal_cell_49_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,19),
			fetch              => s_fetch(49,19),
			data_in            => s_data_in(49,19),
			data_out           => s_data_out(49,19),
			out1               => s_out1(49,19),
			out2               => s_out2(49,19),
			lock_lower_row_out => s_locks_lower_out(49,19),
			lock_lower_row_in  => s_locks_lower_in(49,19),
			in1                => s_in1(49,19),
			in2                => s_in2(49,19),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(19)
		);
	s_in1(49,19)            <= s_out1(50,19);
	s_in2(49,19)            <= s_out2(50,20);
	s_locks_lower_in(49,19) <= s_locks_lower_out(50,19);

		normal_cell_49_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,20),
			fetch              => s_fetch(49,20),
			data_in            => s_data_in(49,20),
			data_out           => s_data_out(49,20),
			out1               => s_out1(49,20),
			out2               => s_out2(49,20),
			lock_lower_row_out => s_locks_lower_out(49,20),
			lock_lower_row_in  => s_locks_lower_in(49,20),
			in1                => s_in1(49,20),
			in2                => s_in2(49,20),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(20)
		);
	s_in1(49,20)            <= s_out1(50,20);
	s_in2(49,20)            <= s_out2(50,21);
	s_locks_lower_in(49,20) <= s_locks_lower_out(50,20);

		normal_cell_49_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,21),
			fetch              => s_fetch(49,21),
			data_in            => s_data_in(49,21),
			data_out           => s_data_out(49,21),
			out1               => s_out1(49,21),
			out2               => s_out2(49,21),
			lock_lower_row_out => s_locks_lower_out(49,21),
			lock_lower_row_in  => s_locks_lower_in(49,21),
			in1                => s_in1(49,21),
			in2                => s_in2(49,21),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(21)
		);
	s_in1(49,21)            <= s_out1(50,21);
	s_in2(49,21)            <= s_out2(50,22);
	s_locks_lower_in(49,21) <= s_locks_lower_out(50,21);

		normal_cell_49_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,22),
			fetch              => s_fetch(49,22),
			data_in            => s_data_in(49,22),
			data_out           => s_data_out(49,22),
			out1               => s_out1(49,22),
			out2               => s_out2(49,22),
			lock_lower_row_out => s_locks_lower_out(49,22),
			lock_lower_row_in  => s_locks_lower_in(49,22),
			in1                => s_in1(49,22),
			in2                => s_in2(49,22),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(22)
		);
	s_in1(49,22)            <= s_out1(50,22);
	s_in2(49,22)            <= s_out2(50,23);
	s_locks_lower_in(49,22) <= s_locks_lower_out(50,22);

		normal_cell_49_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,23),
			fetch              => s_fetch(49,23),
			data_in            => s_data_in(49,23),
			data_out           => s_data_out(49,23),
			out1               => s_out1(49,23),
			out2               => s_out2(49,23),
			lock_lower_row_out => s_locks_lower_out(49,23),
			lock_lower_row_in  => s_locks_lower_in(49,23),
			in1                => s_in1(49,23),
			in2                => s_in2(49,23),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(23)
		);
	s_in1(49,23)            <= s_out1(50,23);
	s_in2(49,23)            <= s_out2(50,24);
	s_locks_lower_in(49,23) <= s_locks_lower_out(50,23);

		normal_cell_49_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,24),
			fetch              => s_fetch(49,24),
			data_in            => s_data_in(49,24),
			data_out           => s_data_out(49,24),
			out1               => s_out1(49,24),
			out2               => s_out2(49,24),
			lock_lower_row_out => s_locks_lower_out(49,24),
			lock_lower_row_in  => s_locks_lower_in(49,24),
			in1                => s_in1(49,24),
			in2                => s_in2(49,24),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(24)
		);
	s_in1(49,24)            <= s_out1(50,24);
	s_in2(49,24)            <= s_out2(50,25);
	s_locks_lower_in(49,24) <= s_locks_lower_out(50,24);

		normal_cell_49_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,25),
			fetch              => s_fetch(49,25),
			data_in            => s_data_in(49,25),
			data_out           => s_data_out(49,25),
			out1               => s_out1(49,25),
			out2               => s_out2(49,25),
			lock_lower_row_out => s_locks_lower_out(49,25),
			lock_lower_row_in  => s_locks_lower_in(49,25),
			in1                => s_in1(49,25),
			in2                => s_in2(49,25),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(25)
		);
	s_in1(49,25)            <= s_out1(50,25);
	s_in2(49,25)            <= s_out2(50,26);
	s_locks_lower_in(49,25) <= s_locks_lower_out(50,25);

		normal_cell_49_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,26),
			fetch              => s_fetch(49,26),
			data_in            => s_data_in(49,26),
			data_out           => s_data_out(49,26),
			out1               => s_out1(49,26),
			out2               => s_out2(49,26),
			lock_lower_row_out => s_locks_lower_out(49,26),
			lock_lower_row_in  => s_locks_lower_in(49,26),
			in1                => s_in1(49,26),
			in2                => s_in2(49,26),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(26)
		);
	s_in1(49,26)            <= s_out1(50,26);
	s_in2(49,26)            <= s_out2(50,27);
	s_locks_lower_in(49,26) <= s_locks_lower_out(50,26);

		normal_cell_49_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,27),
			fetch              => s_fetch(49,27),
			data_in            => s_data_in(49,27),
			data_out           => s_data_out(49,27),
			out1               => s_out1(49,27),
			out2               => s_out2(49,27),
			lock_lower_row_out => s_locks_lower_out(49,27),
			lock_lower_row_in  => s_locks_lower_in(49,27),
			in1                => s_in1(49,27),
			in2                => s_in2(49,27),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(27)
		);
	s_in1(49,27)            <= s_out1(50,27);
	s_in2(49,27)            <= s_out2(50,28);
	s_locks_lower_in(49,27) <= s_locks_lower_out(50,27);

		normal_cell_49_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,28),
			fetch              => s_fetch(49,28),
			data_in            => s_data_in(49,28),
			data_out           => s_data_out(49,28),
			out1               => s_out1(49,28),
			out2               => s_out2(49,28),
			lock_lower_row_out => s_locks_lower_out(49,28),
			lock_lower_row_in  => s_locks_lower_in(49,28),
			in1                => s_in1(49,28),
			in2                => s_in2(49,28),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(28)
		);
	s_in1(49,28)            <= s_out1(50,28);
	s_in2(49,28)            <= s_out2(50,29);
	s_locks_lower_in(49,28) <= s_locks_lower_out(50,28);

		normal_cell_49_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,29),
			fetch              => s_fetch(49,29),
			data_in            => s_data_in(49,29),
			data_out           => s_data_out(49,29),
			out1               => s_out1(49,29),
			out2               => s_out2(49,29),
			lock_lower_row_out => s_locks_lower_out(49,29),
			lock_lower_row_in  => s_locks_lower_in(49,29),
			in1                => s_in1(49,29),
			in2                => s_in2(49,29),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(29)
		);
	s_in1(49,29)            <= s_out1(50,29);
	s_in2(49,29)            <= s_out2(50,30);
	s_locks_lower_in(49,29) <= s_locks_lower_out(50,29);

		normal_cell_49_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,30),
			fetch              => s_fetch(49,30),
			data_in            => s_data_in(49,30),
			data_out           => s_data_out(49,30),
			out1               => s_out1(49,30),
			out2               => s_out2(49,30),
			lock_lower_row_out => s_locks_lower_out(49,30),
			lock_lower_row_in  => s_locks_lower_in(49,30),
			in1                => s_in1(49,30),
			in2                => s_in2(49,30),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(30)
		);
	s_in1(49,30)            <= s_out1(50,30);
	s_in2(49,30)            <= s_out2(50,31);
	s_locks_lower_in(49,30) <= s_locks_lower_out(50,30);

		normal_cell_49_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,31),
			fetch              => s_fetch(49,31),
			data_in            => s_data_in(49,31),
			data_out           => s_data_out(49,31),
			out1               => s_out1(49,31),
			out2               => s_out2(49,31),
			lock_lower_row_out => s_locks_lower_out(49,31),
			lock_lower_row_in  => s_locks_lower_in(49,31),
			in1                => s_in1(49,31),
			in2                => s_in2(49,31),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(31)
		);
	s_in1(49,31)            <= s_out1(50,31);
	s_in2(49,31)            <= s_out2(50,32);
	s_locks_lower_in(49,31) <= s_locks_lower_out(50,31);

		normal_cell_49_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,32),
			fetch              => s_fetch(49,32),
			data_in            => s_data_in(49,32),
			data_out           => s_data_out(49,32),
			out1               => s_out1(49,32),
			out2               => s_out2(49,32),
			lock_lower_row_out => s_locks_lower_out(49,32),
			lock_lower_row_in  => s_locks_lower_in(49,32),
			in1                => s_in1(49,32),
			in2                => s_in2(49,32),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(32)
		);
	s_in1(49,32)            <= s_out1(50,32);
	s_in2(49,32)            <= s_out2(50,33);
	s_locks_lower_in(49,32) <= s_locks_lower_out(50,32);

		normal_cell_49_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,33),
			fetch              => s_fetch(49,33),
			data_in            => s_data_in(49,33),
			data_out           => s_data_out(49,33),
			out1               => s_out1(49,33),
			out2               => s_out2(49,33),
			lock_lower_row_out => s_locks_lower_out(49,33),
			lock_lower_row_in  => s_locks_lower_in(49,33),
			in1                => s_in1(49,33),
			in2                => s_in2(49,33),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(33)
		);
	s_in1(49,33)            <= s_out1(50,33);
	s_in2(49,33)            <= s_out2(50,34);
	s_locks_lower_in(49,33) <= s_locks_lower_out(50,33);

		normal_cell_49_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,34),
			fetch              => s_fetch(49,34),
			data_in            => s_data_in(49,34),
			data_out           => s_data_out(49,34),
			out1               => s_out1(49,34),
			out2               => s_out2(49,34),
			lock_lower_row_out => s_locks_lower_out(49,34),
			lock_lower_row_in  => s_locks_lower_in(49,34),
			in1                => s_in1(49,34),
			in2                => s_in2(49,34),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(34)
		);
	s_in1(49,34)            <= s_out1(50,34);
	s_in2(49,34)            <= s_out2(50,35);
	s_locks_lower_in(49,34) <= s_locks_lower_out(50,34);

		normal_cell_49_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,35),
			fetch              => s_fetch(49,35),
			data_in            => s_data_in(49,35),
			data_out           => s_data_out(49,35),
			out1               => s_out1(49,35),
			out2               => s_out2(49,35),
			lock_lower_row_out => s_locks_lower_out(49,35),
			lock_lower_row_in  => s_locks_lower_in(49,35),
			in1                => s_in1(49,35),
			in2                => s_in2(49,35),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(35)
		);
	s_in1(49,35)            <= s_out1(50,35);
	s_in2(49,35)            <= s_out2(50,36);
	s_locks_lower_in(49,35) <= s_locks_lower_out(50,35);

		normal_cell_49_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,36),
			fetch              => s_fetch(49,36),
			data_in            => s_data_in(49,36),
			data_out           => s_data_out(49,36),
			out1               => s_out1(49,36),
			out2               => s_out2(49,36),
			lock_lower_row_out => s_locks_lower_out(49,36),
			lock_lower_row_in  => s_locks_lower_in(49,36),
			in1                => s_in1(49,36),
			in2                => s_in2(49,36),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(36)
		);
	s_in1(49,36)            <= s_out1(50,36);
	s_in2(49,36)            <= s_out2(50,37);
	s_locks_lower_in(49,36) <= s_locks_lower_out(50,36);

		normal_cell_49_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,37),
			fetch              => s_fetch(49,37),
			data_in            => s_data_in(49,37),
			data_out           => s_data_out(49,37),
			out1               => s_out1(49,37),
			out2               => s_out2(49,37),
			lock_lower_row_out => s_locks_lower_out(49,37),
			lock_lower_row_in  => s_locks_lower_in(49,37),
			in1                => s_in1(49,37),
			in2                => s_in2(49,37),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(37)
		);
	s_in1(49,37)            <= s_out1(50,37);
	s_in2(49,37)            <= s_out2(50,38);
	s_locks_lower_in(49,37) <= s_locks_lower_out(50,37);

		normal_cell_49_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,38),
			fetch              => s_fetch(49,38),
			data_in            => s_data_in(49,38),
			data_out           => s_data_out(49,38),
			out1               => s_out1(49,38),
			out2               => s_out2(49,38),
			lock_lower_row_out => s_locks_lower_out(49,38),
			lock_lower_row_in  => s_locks_lower_in(49,38),
			in1                => s_in1(49,38),
			in2                => s_in2(49,38),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(38)
		);
	s_in1(49,38)            <= s_out1(50,38);
	s_in2(49,38)            <= s_out2(50,39);
	s_locks_lower_in(49,38) <= s_locks_lower_out(50,38);

		normal_cell_49_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,39),
			fetch              => s_fetch(49,39),
			data_in            => s_data_in(49,39),
			data_out           => s_data_out(49,39),
			out1               => s_out1(49,39),
			out2               => s_out2(49,39),
			lock_lower_row_out => s_locks_lower_out(49,39),
			lock_lower_row_in  => s_locks_lower_in(49,39),
			in1                => s_in1(49,39),
			in2                => s_in2(49,39),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(39)
		);
	s_in1(49,39)            <= s_out1(50,39);
	s_in2(49,39)            <= s_out2(50,40);
	s_locks_lower_in(49,39) <= s_locks_lower_out(50,39);

		normal_cell_49_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,40),
			fetch              => s_fetch(49,40),
			data_in            => s_data_in(49,40),
			data_out           => s_data_out(49,40),
			out1               => s_out1(49,40),
			out2               => s_out2(49,40),
			lock_lower_row_out => s_locks_lower_out(49,40),
			lock_lower_row_in  => s_locks_lower_in(49,40),
			in1                => s_in1(49,40),
			in2                => s_in2(49,40),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(40)
		);
	s_in1(49,40)            <= s_out1(50,40);
	s_in2(49,40)            <= s_out2(50,41);
	s_locks_lower_in(49,40) <= s_locks_lower_out(50,40);

		normal_cell_49_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,41),
			fetch              => s_fetch(49,41),
			data_in            => s_data_in(49,41),
			data_out           => s_data_out(49,41),
			out1               => s_out1(49,41),
			out2               => s_out2(49,41),
			lock_lower_row_out => s_locks_lower_out(49,41),
			lock_lower_row_in  => s_locks_lower_in(49,41),
			in1                => s_in1(49,41),
			in2                => s_in2(49,41),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(41)
		);
	s_in1(49,41)            <= s_out1(50,41);
	s_in2(49,41)            <= s_out2(50,42);
	s_locks_lower_in(49,41) <= s_locks_lower_out(50,41);

		normal_cell_49_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,42),
			fetch              => s_fetch(49,42),
			data_in            => s_data_in(49,42),
			data_out           => s_data_out(49,42),
			out1               => s_out1(49,42),
			out2               => s_out2(49,42),
			lock_lower_row_out => s_locks_lower_out(49,42),
			lock_lower_row_in  => s_locks_lower_in(49,42),
			in1                => s_in1(49,42),
			in2                => s_in2(49,42),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(42)
		);
	s_in1(49,42)            <= s_out1(50,42);
	s_in2(49,42)            <= s_out2(50,43);
	s_locks_lower_in(49,42) <= s_locks_lower_out(50,42);

		normal_cell_49_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,43),
			fetch              => s_fetch(49,43),
			data_in            => s_data_in(49,43),
			data_out           => s_data_out(49,43),
			out1               => s_out1(49,43),
			out2               => s_out2(49,43),
			lock_lower_row_out => s_locks_lower_out(49,43),
			lock_lower_row_in  => s_locks_lower_in(49,43),
			in1                => s_in1(49,43),
			in2                => s_in2(49,43),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(43)
		);
	s_in1(49,43)            <= s_out1(50,43);
	s_in2(49,43)            <= s_out2(50,44);
	s_locks_lower_in(49,43) <= s_locks_lower_out(50,43);

		normal_cell_49_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,44),
			fetch              => s_fetch(49,44),
			data_in            => s_data_in(49,44),
			data_out           => s_data_out(49,44),
			out1               => s_out1(49,44),
			out2               => s_out2(49,44),
			lock_lower_row_out => s_locks_lower_out(49,44),
			lock_lower_row_in  => s_locks_lower_in(49,44),
			in1                => s_in1(49,44),
			in2                => s_in2(49,44),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(44)
		);
	s_in1(49,44)            <= s_out1(50,44);
	s_in2(49,44)            <= s_out2(50,45);
	s_locks_lower_in(49,44) <= s_locks_lower_out(50,44);

		normal_cell_49_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,45),
			fetch              => s_fetch(49,45),
			data_in            => s_data_in(49,45),
			data_out           => s_data_out(49,45),
			out1               => s_out1(49,45),
			out2               => s_out2(49,45),
			lock_lower_row_out => s_locks_lower_out(49,45),
			lock_lower_row_in  => s_locks_lower_in(49,45),
			in1                => s_in1(49,45),
			in2                => s_in2(49,45),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(45)
		);
	s_in1(49,45)            <= s_out1(50,45);
	s_in2(49,45)            <= s_out2(50,46);
	s_locks_lower_in(49,45) <= s_locks_lower_out(50,45);

		normal_cell_49_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,46),
			fetch              => s_fetch(49,46),
			data_in            => s_data_in(49,46),
			data_out           => s_data_out(49,46),
			out1               => s_out1(49,46),
			out2               => s_out2(49,46),
			lock_lower_row_out => s_locks_lower_out(49,46),
			lock_lower_row_in  => s_locks_lower_in(49,46),
			in1                => s_in1(49,46),
			in2                => s_in2(49,46),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(46)
		);
	s_in1(49,46)            <= s_out1(50,46);
	s_in2(49,46)            <= s_out2(50,47);
	s_locks_lower_in(49,46) <= s_locks_lower_out(50,46);

		normal_cell_49_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,47),
			fetch              => s_fetch(49,47),
			data_in            => s_data_in(49,47),
			data_out           => s_data_out(49,47),
			out1               => s_out1(49,47),
			out2               => s_out2(49,47),
			lock_lower_row_out => s_locks_lower_out(49,47),
			lock_lower_row_in  => s_locks_lower_in(49,47),
			in1                => s_in1(49,47),
			in2                => s_in2(49,47),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(47)
		);
	s_in1(49,47)            <= s_out1(50,47);
	s_in2(49,47)            <= s_out2(50,48);
	s_locks_lower_in(49,47) <= s_locks_lower_out(50,47);

		normal_cell_49_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,48),
			fetch              => s_fetch(49,48),
			data_in            => s_data_in(49,48),
			data_out           => s_data_out(49,48),
			out1               => s_out1(49,48),
			out2               => s_out2(49,48),
			lock_lower_row_out => s_locks_lower_out(49,48),
			lock_lower_row_in  => s_locks_lower_in(49,48),
			in1                => s_in1(49,48),
			in2                => s_in2(49,48),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(48)
		);
	s_in1(49,48)            <= s_out1(50,48);
	s_in2(49,48)            <= s_out2(50,49);
	s_locks_lower_in(49,48) <= s_locks_lower_out(50,48);

		normal_cell_49_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,49),
			fetch              => s_fetch(49,49),
			data_in            => s_data_in(49,49),
			data_out           => s_data_out(49,49),
			out1               => s_out1(49,49),
			out2               => s_out2(49,49),
			lock_lower_row_out => s_locks_lower_out(49,49),
			lock_lower_row_in  => s_locks_lower_in(49,49),
			in1                => s_in1(49,49),
			in2                => s_in2(49,49),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(49)
		);
	s_in1(49,49)            <= s_out1(50,49);
	s_in2(49,49)            <= s_out2(50,50);
	s_locks_lower_in(49,49) <= s_locks_lower_out(50,49);

		normal_cell_49_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,50),
			fetch              => s_fetch(49,50),
			data_in            => s_data_in(49,50),
			data_out           => s_data_out(49,50),
			out1               => s_out1(49,50),
			out2               => s_out2(49,50),
			lock_lower_row_out => s_locks_lower_out(49,50),
			lock_lower_row_in  => s_locks_lower_in(49,50),
			in1                => s_in1(49,50),
			in2                => s_in2(49,50),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(50)
		);
	s_in1(49,50)            <= s_out1(50,50);
	s_in2(49,50)            <= s_out2(50,51);
	s_locks_lower_in(49,50) <= s_locks_lower_out(50,50);

		normal_cell_49_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,51),
			fetch              => s_fetch(49,51),
			data_in            => s_data_in(49,51),
			data_out           => s_data_out(49,51),
			out1               => s_out1(49,51),
			out2               => s_out2(49,51),
			lock_lower_row_out => s_locks_lower_out(49,51),
			lock_lower_row_in  => s_locks_lower_in(49,51),
			in1                => s_in1(49,51),
			in2                => s_in2(49,51),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(51)
		);
	s_in1(49,51)            <= s_out1(50,51);
	s_in2(49,51)            <= s_out2(50,52);
	s_locks_lower_in(49,51) <= s_locks_lower_out(50,51);

		normal_cell_49_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,52),
			fetch              => s_fetch(49,52),
			data_in            => s_data_in(49,52),
			data_out           => s_data_out(49,52),
			out1               => s_out1(49,52),
			out2               => s_out2(49,52),
			lock_lower_row_out => s_locks_lower_out(49,52),
			lock_lower_row_in  => s_locks_lower_in(49,52),
			in1                => s_in1(49,52),
			in2                => s_in2(49,52),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(52)
		);
	s_in1(49,52)            <= s_out1(50,52);
	s_in2(49,52)            <= s_out2(50,53);
	s_locks_lower_in(49,52) <= s_locks_lower_out(50,52);

		normal_cell_49_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,53),
			fetch              => s_fetch(49,53),
			data_in            => s_data_in(49,53),
			data_out           => s_data_out(49,53),
			out1               => s_out1(49,53),
			out2               => s_out2(49,53),
			lock_lower_row_out => s_locks_lower_out(49,53),
			lock_lower_row_in  => s_locks_lower_in(49,53),
			in1                => s_in1(49,53),
			in2                => s_in2(49,53),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(53)
		);
	s_in1(49,53)            <= s_out1(50,53);
	s_in2(49,53)            <= s_out2(50,54);
	s_locks_lower_in(49,53) <= s_locks_lower_out(50,53);

		normal_cell_49_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,54),
			fetch              => s_fetch(49,54),
			data_in            => s_data_in(49,54),
			data_out           => s_data_out(49,54),
			out1               => s_out1(49,54),
			out2               => s_out2(49,54),
			lock_lower_row_out => s_locks_lower_out(49,54),
			lock_lower_row_in  => s_locks_lower_in(49,54),
			in1                => s_in1(49,54),
			in2                => s_in2(49,54),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(54)
		);
	s_in1(49,54)            <= s_out1(50,54);
	s_in2(49,54)            <= s_out2(50,55);
	s_locks_lower_in(49,54) <= s_locks_lower_out(50,54);

		normal_cell_49_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,55),
			fetch              => s_fetch(49,55),
			data_in            => s_data_in(49,55),
			data_out           => s_data_out(49,55),
			out1               => s_out1(49,55),
			out2               => s_out2(49,55),
			lock_lower_row_out => s_locks_lower_out(49,55),
			lock_lower_row_in  => s_locks_lower_in(49,55),
			in1                => s_in1(49,55),
			in2                => s_in2(49,55),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(55)
		);
	s_in1(49,55)            <= s_out1(50,55);
	s_in2(49,55)            <= s_out2(50,56);
	s_locks_lower_in(49,55) <= s_locks_lower_out(50,55);

		normal_cell_49_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,56),
			fetch              => s_fetch(49,56),
			data_in            => s_data_in(49,56),
			data_out           => s_data_out(49,56),
			out1               => s_out1(49,56),
			out2               => s_out2(49,56),
			lock_lower_row_out => s_locks_lower_out(49,56),
			lock_lower_row_in  => s_locks_lower_in(49,56),
			in1                => s_in1(49,56),
			in2                => s_in2(49,56),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(56)
		);
	s_in1(49,56)            <= s_out1(50,56);
	s_in2(49,56)            <= s_out2(50,57);
	s_locks_lower_in(49,56) <= s_locks_lower_out(50,56);

		normal_cell_49_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,57),
			fetch              => s_fetch(49,57),
			data_in            => s_data_in(49,57),
			data_out           => s_data_out(49,57),
			out1               => s_out1(49,57),
			out2               => s_out2(49,57),
			lock_lower_row_out => s_locks_lower_out(49,57),
			lock_lower_row_in  => s_locks_lower_in(49,57),
			in1                => s_in1(49,57),
			in2                => s_in2(49,57),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(57)
		);
	s_in1(49,57)            <= s_out1(50,57);
	s_in2(49,57)            <= s_out2(50,58);
	s_locks_lower_in(49,57) <= s_locks_lower_out(50,57);

		normal_cell_49_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,58),
			fetch              => s_fetch(49,58),
			data_in            => s_data_in(49,58),
			data_out           => s_data_out(49,58),
			out1               => s_out1(49,58),
			out2               => s_out2(49,58),
			lock_lower_row_out => s_locks_lower_out(49,58),
			lock_lower_row_in  => s_locks_lower_in(49,58),
			in1                => s_in1(49,58),
			in2                => s_in2(49,58),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(58)
		);
	s_in1(49,58)            <= s_out1(50,58);
	s_in2(49,58)            <= s_out2(50,59);
	s_locks_lower_in(49,58) <= s_locks_lower_out(50,58);

		normal_cell_49_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,59),
			fetch              => s_fetch(49,59),
			data_in            => s_data_in(49,59),
			data_out           => s_data_out(49,59),
			out1               => s_out1(49,59),
			out2               => s_out2(49,59),
			lock_lower_row_out => s_locks_lower_out(49,59),
			lock_lower_row_in  => s_locks_lower_in(49,59),
			in1                => s_in1(49,59),
			in2                => s_in2(49,59),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(59)
		);
	s_in1(49,59)            <= s_out1(50,59);
	s_in2(49,59)            <= s_out2(50,60);
	s_locks_lower_in(49,59) <= s_locks_lower_out(50,59);

		last_col_cell_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(49,60),
			fetch              => s_fetch(49,60),
			data_in            => s_data_in(49,60),
			data_out           => s_data_out(49,60),
			out1               => s_out1(49,60),
			out2               => s_out2(49,60),
			lock_lower_row_out => s_locks_lower_out(49,60),
			lock_lower_row_in  => s_locks_lower_in(49,60),
			in1                => s_in1(49,60),
			in2                => (others => '0'),
			lock_row           => s_locks(49),
			piv_found          => s_piv_found,
			row_data           => s_row_data(49),
			col_data           => s_col_data(60)
		);
	s_in1(49,60)            <= s_out1(50,60);
	s_locks_lower_in(49,60) <= s_locks_lower_out(50,60);

		normal_cell_50_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,1),
			fetch              => s_fetch(50,1),
			data_in            => s_data_in(50,1),
			data_out           => s_data_out(50,1),
			out1               => s_out1(50,1),
			out2               => s_out2(50,1),
			lock_lower_row_out => s_locks_lower_out(50,1),
			lock_lower_row_in  => s_locks_lower_in(50,1),
			in1                => s_in1(50,1),
			in2                => s_in2(50,1),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(1)
		);
	s_in1(50,1)            <= s_out1(51,1);
	s_in2(50,1)            <= s_out2(51,2);
	s_locks_lower_in(50,1) <= s_locks_lower_out(51,1);

		normal_cell_50_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,2),
			fetch              => s_fetch(50,2),
			data_in            => s_data_in(50,2),
			data_out           => s_data_out(50,2),
			out1               => s_out1(50,2),
			out2               => s_out2(50,2),
			lock_lower_row_out => s_locks_lower_out(50,2),
			lock_lower_row_in  => s_locks_lower_in(50,2),
			in1                => s_in1(50,2),
			in2                => s_in2(50,2),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(2)
		);
	s_in1(50,2)            <= s_out1(51,2);
	s_in2(50,2)            <= s_out2(51,3);
	s_locks_lower_in(50,2) <= s_locks_lower_out(51,2);

		normal_cell_50_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,3),
			fetch              => s_fetch(50,3),
			data_in            => s_data_in(50,3),
			data_out           => s_data_out(50,3),
			out1               => s_out1(50,3),
			out2               => s_out2(50,3),
			lock_lower_row_out => s_locks_lower_out(50,3),
			lock_lower_row_in  => s_locks_lower_in(50,3),
			in1                => s_in1(50,3),
			in2                => s_in2(50,3),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(3)
		);
	s_in1(50,3)            <= s_out1(51,3);
	s_in2(50,3)            <= s_out2(51,4);
	s_locks_lower_in(50,3) <= s_locks_lower_out(51,3);

		normal_cell_50_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,4),
			fetch              => s_fetch(50,4),
			data_in            => s_data_in(50,4),
			data_out           => s_data_out(50,4),
			out1               => s_out1(50,4),
			out2               => s_out2(50,4),
			lock_lower_row_out => s_locks_lower_out(50,4),
			lock_lower_row_in  => s_locks_lower_in(50,4),
			in1                => s_in1(50,4),
			in2                => s_in2(50,4),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(4)
		);
	s_in1(50,4)            <= s_out1(51,4);
	s_in2(50,4)            <= s_out2(51,5);
	s_locks_lower_in(50,4) <= s_locks_lower_out(51,4);

		normal_cell_50_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,5),
			fetch              => s_fetch(50,5),
			data_in            => s_data_in(50,5),
			data_out           => s_data_out(50,5),
			out1               => s_out1(50,5),
			out2               => s_out2(50,5),
			lock_lower_row_out => s_locks_lower_out(50,5),
			lock_lower_row_in  => s_locks_lower_in(50,5),
			in1                => s_in1(50,5),
			in2                => s_in2(50,5),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(5)
		);
	s_in1(50,5)            <= s_out1(51,5);
	s_in2(50,5)            <= s_out2(51,6);
	s_locks_lower_in(50,5) <= s_locks_lower_out(51,5);

		normal_cell_50_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,6),
			fetch              => s_fetch(50,6),
			data_in            => s_data_in(50,6),
			data_out           => s_data_out(50,6),
			out1               => s_out1(50,6),
			out2               => s_out2(50,6),
			lock_lower_row_out => s_locks_lower_out(50,6),
			lock_lower_row_in  => s_locks_lower_in(50,6),
			in1                => s_in1(50,6),
			in2                => s_in2(50,6),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(6)
		);
	s_in1(50,6)            <= s_out1(51,6);
	s_in2(50,6)            <= s_out2(51,7);
	s_locks_lower_in(50,6) <= s_locks_lower_out(51,6);

		normal_cell_50_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,7),
			fetch              => s_fetch(50,7),
			data_in            => s_data_in(50,7),
			data_out           => s_data_out(50,7),
			out1               => s_out1(50,7),
			out2               => s_out2(50,7),
			lock_lower_row_out => s_locks_lower_out(50,7),
			lock_lower_row_in  => s_locks_lower_in(50,7),
			in1                => s_in1(50,7),
			in2                => s_in2(50,7),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(7)
		);
	s_in1(50,7)            <= s_out1(51,7);
	s_in2(50,7)            <= s_out2(51,8);
	s_locks_lower_in(50,7) <= s_locks_lower_out(51,7);

		normal_cell_50_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,8),
			fetch              => s_fetch(50,8),
			data_in            => s_data_in(50,8),
			data_out           => s_data_out(50,8),
			out1               => s_out1(50,8),
			out2               => s_out2(50,8),
			lock_lower_row_out => s_locks_lower_out(50,8),
			lock_lower_row_in  => s_locks_lower_in(50,8),
			in1                => s_in1(50,8),
			in2                => s_in2(50,8),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(8)
		);
	s_in1(50,8)            <= s_out1(51,8);
	s_in2(50,8)            <= s_out2(51,9);
	s_locks_lower_in(50,8) <= s_locks_lower_out(51,8);

		normal_cell_50_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,9),
			fetch              => s_fetch(50,9),
			data_in            => s_data_in(50,9),
			data_out           => s_data_out(50,9),
			out1               => s_out1(50,9),
			out2               => s_out2(50,9),
			lock_lower_row_out => s_locks_lower_out(50,9),
			lock_lower_row_in  => s_locks_lower_in(50,9),
			in1                => s_in1(50,9),
			in2                => s_in2(50,9),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(9)
		);
	s_in1(50,9)            <= s_out1(51,9);
	s_in2(50,9)            <= s_out2(51,10);
	s_locks_lower_in(50,9) <= s_locks_lower_out(51,9);

		normal_cell_50_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,10),
			fetch              => s_fetch(50,10),
			data_in            => s_data_in(50,10),
			data_out           => s_data_out(50,10),
			out1               => s_out1(50,10),
			out2               => s_out2(50,10),
			lock_lower_row_out => s_locks_lower_out(50,10),
			lock_lower_row_in  => s_locks_lower_in(50,10),
			in1                => s_in1(50,10),
			in2                => s_in2(50,10),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(10)
		);
	s_in1(50,10)            <= s_out1(51,10);
	s_in2(50,10)            <= s_out2(51,11);
	s_locks_lower_in(50,10) <= s_locks_lower_out(51,10);

		normal_cell_50_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,11),
			fetch              => s_fetch(50,11),
			data_in            => s_data_in(50,11),
			data_out           => s_data_out(50,11),
			out1               => s_out1(50,11),
			out2               => s_out2(50,11),
			lock_lower_row_out => s_locks_lower_out(50,11),
			lock_lower_row_in  => s_locks_lower_in(50,11),
			in1                => s_in1(50,11),
			in2                => s_in2(50,11),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(11)
		);
	s_in1(50,11)            <= s_out1(51,11);
	s_in2(50,11)            <= s_out2(51,12);
	s_locks_lower_in(50,11) <= s_locks_lower_out(51,11);

		normal_cell_50_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,12),
			fetch              => s_fetch(50,12),
			data_in            => s_data_in(50,12),
			data_out           => s_data_out(50,12),
			out1               => s_out1(50,12),
			out2               => s_out2(50,12),
			lock_lower_row_out => s_locks_lower_out(50,12),
			lock_lower_row_in  => s_locks_lower_in(50,12),
			in1                => s_in1(50,12),
			in2                => s_in2(50,12),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(12)
		);
	s_in1(50,12)            <= s_out1(51,12);
	s_in2(50,12)            <= s_out2(51,13);
	s_locks_lower_in(50,12) <= s_locks_lower_out(51,12);

		normal_cell_50_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,13),
			fetch              => s_fetch(50,13),
			data_in            => s_data_in(50,13),
			data_out           => s_data_out(50,13),
			out1               => s_out1(50,13),
			out2               => s_out2(50,13),
			lock_lower_row_out => s_locks_lower_out(50,13),
			lock_lower_row_in  => s_locks_lower_in(50,13),
			in1                => s_in1(50,13),
			in2                => s_in2(50,13),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(13)
		);
	s_in1(50,13)            <= s_out1(51,13);
	s_in2(50,13)            <= s_out2(51,14);
	s_locks_lower_in(50,13) <= s_locks_lower_out(51,13);

		normal_cell_50_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,14),
			fetch              => s_fetch(50,14),
			data_in            => s_data_in(50,14),
			data_out           => s_data_out(50,14),
			out1               => s_out1(50,14),
			out2               => s_out2(50,14),
			lock_lower_row_out => s_locks_lower_out(50,14),
			lock_lower_row_in  => s_locks_lower_in(50,14),
			in1                => s_in1(50,14),
			in2                => s_in2(50,14),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(14)
		);
	s_in1(50,14)            <= s_out1(51,14);
	s_in2(50,14)            <= s_out2(51,15);
	s_locks_lower_in(50,14) <= s_locks_lower_out(51,14);

		normal_cell_50_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,15),
			fetch              => s_fetch(50,15),
			data_in            => s_data_in(50,15),
			data_out           => s_data_out(50,15),
			out1               => s_out1(50,15),
			out2               => s_out2(50,15),
			lock_lower_row_out => s_locks_lower_out(50,15),
			lock_lower_row_in  => s_locks_lower_in(50,15),
			in1                => s_in1(50,15),
			in2                => s_in2(50,15),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(15)
		);
	s_in1(50,15)            <= s_out1(51,15);
	s_in2(50,15)            <= s_out2(51,16);
	s_locks_lower_in(50,15) <= s_locks_lower_out(51,15);

		normal_cell_50_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,16),
			fetch              => s_fetch(50,16),
			data_in            => s_data_in(50,16),
			data_out           => s_data_out(50,16),
			out1               => s_out1(50,16),
			out2               => s_out2(50,16),
			lock_lower_row_out => s_locks_lower_out(50,16),
			lock_lower_row_in  => s_locks_lower_in(50,16),
			in1                => s_in1(50,16),
			in2                => s_in2(50,16),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(16)
		);
	s_in1(50,16)            <= s_out1(51,16);
	s_in2(50,16)            <= s_out2(51,17);
	s_locks_lower_in(50,16) <= s_locks_lower_out(51,16);

		normal_cell_50_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,17),
			fetch              => s_fetch(50,17),
			data_in            => s_data_in(50,17),
			data_out           => s_data_out(50,17),
			out1               => s_out1(50,17),
			out2               => s_out2(50,17),
			lock_lower_row_out => s_locks_lower_out(50,17),
			lock_lower_row_in  => s_locks_lower_in(50,17),
			in1                => s_in1(50,17),
			in2                => s_in2(50,17),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(17)
		);
	s_in1(50,17)            <= s_out1(51,17);
	s_in2(50,17)            <= s_out2(51,18);
	s_locks_lower_in(50,17) <= s_locks_lower_out(51,17);

		normal_cell_50_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,18),
			fetch              => s_fetch(50,18),
			data_in            => s_data_in(50,18),
			data_out           => s_data_out(50,18),
			out1               => s_out1(50,18),
			out2               => s_out2(50,18),
			lock_lower_row_out => s_locks_lower_out(50,18),
			lock_lower_row_in  => s_locks_lower_in(50,18),
			in1                => s_in1(50,18),
			in2                => s_in2(50,18),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(18)
		);
	s_in1(50,18)            <= s_out1(51,18);
	s_in2(50,18)            <= s_out2(51,19);
	s_locks_lower_in(50,18) <= s_locks_lower_out(51,18);

		normal_cell_50_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,19),
			fetch              => s_fetch(50,19),
			data_in            => s_data_in(50,19),
			data_out           => s_data_out(50,19),
			out1               => s_out1(50,19),
			out2               => s_out2(50,19),
			lock_lower_row_out => s_locks_lower_out(50,19),
			lock_lower_row_in  => s_locks_lower_in(50,19),
			in1                => s_in1(50,19),
			in2                => s_in2(50,19),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(19)
		);
	s_in1(50,19)            <= s_out1(51,19);
	s_in2(50,19)            <= s_out2(51,20);
	s_locks_lower_in(50,19) <= s_locks_lower_out(51,19);

		normal_cell_50_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,20),
			fetch              => s_fetch(50,20),
			data_in            => s_data_in(50,20),
			data_out           => s_data_out(50,20),
			out1               => s_out1(50,20),
			out2               => s_out2(50,20),
			lock_lower_row_out => s_locks_lower_out(50,20),
			lock_lower_row_in  => s_locks_lower_in(50,20),
			in1                => s_in1(50,20),
			in2                => s_in2(50,20),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(20)
		);
	s_in1(50,20)            <= s_out1(51,20);
	s_in2(50,20)            <= s_out2(51,21);
	s_locks_lower_in(50,20) <= s_locks_lower_out(51,20);

		normal_cell_50_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,21),
			fetch              => s_fetch(50,21),
			data_in            => s_data_in(50,21),
			data_out           => s_data_out(50,21),
			out1               => s_out1(50,21),
			out2               => s_out2(50,21),
			lock_lower_row_out => s_locks_lower_out(50,21),
			lock_lower_row_in  => s_locks_lower_in(50,21),
			in1                => s_in1(50,21),
			in2                => s_in2(50,21),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(21)
		);
	s_in1(50,21)            <= s_out1(51,21);
	s_in2(50,21)            <= s_out2(51,22);
	s_locks_lower_in(50,21) <= s_locks_lower_out(51,21);

		normal_cell_50_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,22),
			fetch              => s_fetch(50,22),
			data_in            => s_data_in(50,22),
			data_out           => s_data_out(50,22),
			out1               => s_out1(50,22),
			out2               => s_out2(50,22),
			lock_lower_row_out => s_locks_lower_out(50,22),
			lock_lower_row_in  => s_locks_lower_in(50,22),
			in1                => s_in1(50,22),
			in2                => s_in2(50,22),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(22)
		);
	s_in1(50,22)            <= s_out1(51,22);
	s_in2(50,22)            <= s_out2(51,23);
	s_locks_lower_in(50,22) <= s_locks_lower_out(51,22);

		normal_cell_50_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,23),
			fetch              => s_fetch(50,23),
			data_in            => s_data_in(50,23),
			data_out           => s_data_out(50,23),
			out1               => s_out1(50,23),
			out2               => s_out2(50,23),
			lock_lower_row_out => s_locks_lower_out(50,23),
			lock_lower_row_in  => s_locks_lower_in(50,23),
			in1                => s_in1(50,23),
			in2                => s_in2(50,23),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(23)
		);
	s_in1(50,23)            <= s_out1(51,23);
	s_in2(50,23)            <= s_out2(51,24);
	s_locks_lower_in(50,23) <= s_locks_lower_out(51,23);

		normal_cell_50_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,24),
			fetch              => s_fetch(50,24),
			data_in            => s_data_in(50,24),
			data_out           => s_data_out(50,24),
			out1               => s_out1(50,24),
			out2               => s_out2(50,24),
			lock_lower_row_out => s_locks_lower_out(50,24),
			lock_lower_row_in  => s_locks_lower_in(50,24),
			in1                => s_in1(50,24),
			in2                => s_in2(50,24),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(24)
		);
	s_in1(50,24)            <= s_out1(51,24);
	s_in2(50,24)            <= s_out2(51,25);
	s_locks_lower_in(50,24) <= s_locks_lower_out(51,24);

		normal_cell_50_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,25),
			fetch              => s_fetch(50,25),
			data_in            => s_data_in(50,25),
			data_out           => s_data_out(50,25),
			out1               => s_out1(50,25),
			out2               => s_out2(50,25),
			lock_lower_row_out => s_locks_lower_out(50,25),
			lock_lower_row_in  => s_locks_lower_in(50,25),
			in1                => s_in1(50,25),
			in2                => s_in2(50,25),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(25)
		);
	s_in1(50,25)            <= s_out1(51,25);
	s_in2(50,25)            <= s_out2(51,26);
	s_locks_lower_in(50,25) <= s_locks_lower_out(51,25);

		normal_cell_50_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,26),
			fetch              => s_fetch(50,26),
			data_in            => s_data_in(50,26),
			data_out           => s_data_out(50,26),
			out1               => s_out1(50,26),
			out2               => s_out2(50,26),
			lock_lower_row_out => s_locks_lower_out(50,26),
			lock_lower_row_in  => s_locks_lower_in(50,26),
			in1                => s_in1(50,26),
			in2                => s_in2(50,26),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(26)
		);
	s_in1(50,26)            <= s_out1(51,26);
	s_in2(50,26)            <= s_out2(51,27);
	s_locks_lower_in(50,26) <= s_locks_lower_out(51,26);

		normal_cell_50_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,27),
			fetch              => s_fetch(50,27),
			data_in            => s_data_in(50,27),
			data_out           => s_data_out(50,27),
			out1               => s_out1(50,27),
			out2               => s_out2(50,27),
			lock_lower_row_out => s_locks_lower_out(50,27),
			lock_lower_row_in  => s_locks_lower_in(50,27),
			in1                => s_in1(50,27),
			in2                => s_in2(50,27),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(27)
		);
	s_in1(50,27)            <= s_out1(51,27);
	s_in2(50,27)            <= s_out2(51,28);
	s_locks_lower_in(50,27) <= s_locks_lower_out(51,27);

		normal_cell_50_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,28),
			fetch              => s_fetch(50,28),
			data_in            => s_data_in(50,28),
			data_out           => s_data_out(50,28),
			out1               => s_out1(50,28),
			out2               => s_out2(50,28),
			lock_lower_row_out => s_locks_lower_out(50,28),
			lock_lower_row_in  => s_locks_lower_in(50,28),
			in1                => s_in1(50,28),
			in2                => s_in2(50,28),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(28)
		);
	s_in1(50,28)            <= s_out1(51,28);
	s_in2(50,28)            <= s_out2(51,29);
	s_locks_lower_in(50,28) <= s_locks_lower_out(51,28);

		normal_cell_50_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,29),
			fetch              => s_fetch(50,29),
			data_in            => s_data_in(50,29),
			data_out           => s_data_out(50,29),
			out1               => s_out1(50,29),
			out2               => s_out2(50,29),
			lock_lower_row_out => s_locks_lower_out(50,29),
			lock_lower_row_in  => s_locks_lower_in(50,29),
			in1                => s_in1(50,29),
			in2                => s_in2(50,29),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(29)
		);
	s_in1(50,29)            <= s_out1(51,29);
	s_in2(50,29)            <= s_out2(51,30);
	s_locks_lower_in(50,29) <= s_locks_lower_out(51,29);

		normal_cell_50_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,30),
			fetch              => s_fetch(50,30),
			data_in            => s_data_in(50,30),
			data_out           => s_data_out(50,30),
			out1               => s_out1(50,30),
			out2               => s_out2(50,30),
			lock_lower_row_out => s_locks_lower_out(50,30),
			lock_lower_row_in  => s_locks_lower_in(50,30),
			in1                => s_in1(50,30),
			in2                => s_in2(50,30),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(30)
		);
	s_in1(50,30)            <= s_out1(51,30);
	s_in2(50,30)            <= s_out2(51,31);
	s_locks_lower_in(50,30) <= s_locks_lower_out(51,30);

		normal_cell_50_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,31),
			fetch              => s_fetch(50,31),
			data_in            => s_data_in(50,31),
			data_out           => s_data_out(50,31),
			out1               => s_out1(50,31),
			out2               => s_out2(50,31),
			lock_lower_row_out => s_locks_lower_out(50,31),
			lock_lower_row_in  => s_locks_lower_in(50,31),
			in1                => s_in1(50,31),
			in2                => s_in2(50,31),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(31)
		);
	s_in1(50,31)            <= s_out1(51,31);
	s_in2(50,31)            <= s_out2(51,32);
	s_locks_lower_in(50,31) <= s_locks_lower_out(51,31);

		normal_cell_50_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,32),
			fetch              => s_fetch(50,32),
			data_in            => s_data_in(50,32),
			data_out           => s_data_out(50,32),
			out1               => s_out1(50,32),
			out2               => s_out2(50,32),
			lock_lower_row_out => s_locks_lower_out(50,32),
			lock_lower_row_in  => s_locks_lower_in(50,32),
			in1                => s_in1(50,32),
			in2                => s_in2(50,32),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(32)
		);
	s_in1(50,32)            <= s_out1(51,32);
	s_in2(50,32)            <= s_out2(51,33);
	s_locks_lower_in(50,32) <= s_locks_lower_out(51,32);

		normal_cell_50_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,33),
			fetch              => s_fetch(50,33),
			data_in            => s_data_in(50,33),
			data_out           => s_data_out(50,33),
			out1               => s_out1(50,33),
			out2               => s_out2(50,33),
			lock_lower_row_out => s_locks_lower_out(50,33),
			lock_lower_row_in  => s_locks_lower_in(50,33),
			in1                => s_in1(50,33),
			in2                => s_in2(50,33),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(33)
		);
	s_in1(50,33)            <= s_out1(51,33);
	s_in2(50,33)            <= s_out2(51,34);
	s_locks_lower_in(50,33) <= s_locks_lower_out(51,33);

		normal_cell_50_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,34),
			fetch              => s_fetch(50,34),
			data_in            => s_data_in(50,34),
			data_out           => s_data_out(50,34),
			out1               => s_out1(50,34),
			out2               => s_out2(50,34),
			lock_lower_row_out => s_locks_lower_out(50,34),
			lock_lower_row_in  => s_locks_lower_in(50,34),
			in1                => s_in1(50,34),
			in2                => s_in2(50,34),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(34)
		);
	s_in1(50,34)            <= s_out1(51,34);
	s_in2(50,34)            <= s_out2(51,35);
	s_locks_lower_in(50,34) <= s_locks_lower_out(51,34);

		normal_cell_50_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,35),
			fetch              => s_fetch(50,35),
			data_in            => s_data_in(50,35),
			data_out           => s_data_out(50,35),
			out1               => s_out1(50,35),
			out2               => s_out2(50,35),
			lock_lower_row_out => s_locks_lower_out(50,35),
			lock_lower_row_in  => s_locks_lower_in(50,35),
			in1                => s_in1(50,35),
			in2                => s_in2(50,35),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(35)
		);
	s_in1(50,35)            <= s_out1(51,35);
	s_in2(50,35)            <= s_out2(51,36);
	s_locks_lower_in(50,35) <= s_locks_lower_out(51,35);

		normal_cell_50_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,36),
			fetch              => s_fetch(50,36),
			data_in            => s_data_in(50,36),
			data_out           => s_data_out(50,36),
			out1               => s_out1(50,36),
			out2               => s_out2(50,36),
			lock_lower_row_out => s_locks_lower_out(50,36),
			lock_lower_row_in  => s_locks_lower_in(50,36),
			in1                => s_in1(50,36),
			in2                => s_in2(50,36),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(36)
		);
	s_in1(50,36)            <= s_out1(51,36);
	s_in2(50,36)            <= s_out2(51,37);
	s_locks_lower_in(50,36) <= s_locks_lower_out(51,36);

		normal_cell_50_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,37),
			fetch              => s_fetch(50,37),
			data_in            => s_data_in(50,37),
			data_out           => s_data_out(50,37),
			out1               => s_out1(50,37),
			out2               => s_out2(50,37),
			lock_lower_row_out => s_locks_lower_out(50,37),
			lock_lower_row_in  => s_locks_lower_in(50,37),
			in1                => s_in1(50,37),
			in2                => s_in2(50,37),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(37)
		);
	s_in1(50,37)            <= s_out1(51,37);
	s_in2(50,37)            <= s_out2(51,38);
	s_locks_lower_in(50,37) <= s_locks_lower_out(51,37);

		normal_cell_50_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,38),
			fetch              => s_fetch(50,38),
			data_in            => s_data_in(50,38),
			data_out           => s_data_out(50,38),
			out1               => s_out1(50,38),
			out2               => s_out2(50,38),
			lock_lower_row_out => s_locks_lower_out(50,38),
			lock_lower_row_in  => s_locks_lower_in(50,38),
			in1                => s_in1(50,38),
			in2                => s_in2(50,38),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(38)
		);
	s_in1(50,38)            <= s_out1(51,38);
	s_in2(50,38)            <= s_out2(51,39);
	s_locks_lower_in(50,38) <= s_locks_lower_out(51,38);

		normal_cell_50_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,39),
			fetch              => s_fetch(50,39),
			data_in            => s_data_in(50,39),
			data_out           => s_data_out(50,39),
			out1               => s_out1(50,39),
			out2               => s_out2(50,39),
			lock_lower_row_out => s_locks_lower_out(50,39),
			lock_lower_row_in  => s_locks_lower_in(50,39),
			in1                => s_in1(50,39),
			in2                => s_in2(50,39),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(39)
		);
	s_in1(50,39)            <= s_out1(51,39);
	s_in2(50,39)            <= s_out2(51,40);
	s_locks_lower_in(50,39) <= s_locks_lower_out(51,39);

		normal_cell_50_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,40),
			fetch              => s_fetch(50,40),
			data_in            => s_data_in(50,40),
			data_out           => s_data_out(50,40),
			out1               => s_out1(50,40),
			out2               => s_out2(50,40),
			lock_lower_row_out => s_locks_lower_out(50,40),
			lock_lower_row_in  => s_locks_lower_in(50,40),
			in1                => s_in1(50,40),
			in2                => s_in2(50,40),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(40)
		);
	s_in1(50,40)            <= s_out1(51,40);
	s_in2(50,40)            <= s_out2(51,41);
	s_locks_lower_in(50,40) <= s_locks_lower_out(51,40);

		normal_cell_50_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,41),
			fetch              => s_fetch(50,41),
			data_in            => s_data_in(50,41),
			data_out           => s_data_out(50,41),
			out1               => s_out1(50,41),
			out2               => s_out2(50,41),
			lock_lower_row_out => s_locks_lower_out(50,41),
			lock_lower_row_in  => s_locks_lower_in(50,41),
			in1                => s_in1(50,41),
			in2                => s_in2(50,41),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(41)
		);
	s_in1(50,41)            <= s_out1(51,41);
	s_in2(50,41)            <= s_out2(51,42);
	s_locks_lower_in(50,41) <= s_locks_lower_out(51,41);

		normal_cell_50_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,42),
			fetch              => s_fetch(50,42),
			data_in            => s_data_in(50,42),
			data_out           => s_data_out(50,42),
			out1               => s_out1(50,42),
			out2               => s_out2(50,42),
			lock_lower_row_out => s_locks_lower_out(50,42),
			lock_lower_row_in  => s_locks_lower_in(50,42),
			in1                => s_in1(50,42),
			in2                => s_in2(50,42),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(42)
		);
	s_in1(50,42)            <= s_out1(51,42);
	s_in2(50,42)            <= s_out2(51,43);
	s_locks_lower_in(50,42) <= s_locks_lower_out(51,42);

		normal_cell_50_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,43),
			fetch              => s_fetch(50,43),
			data_in            => s_data_in(50,43),
			data_out           => s_data_out(50,43),
			out1               => s_out1(50,43),
			out2               => s_out2(50,43),
			lock_lower_row_out => s_locks_lower_out(50,43),
			lock_lower_row_in  => s_locks_lower_in(50,43),
			in1                => s_in1(50,43),
			in2                => s_in2(50,43),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(43)
		);
	s_in1(50,43)            <= s_out1(51,43);
	s_in2(50,43)            <= s_out2(51,44);
	s_locks_lower_in(50,43) <= s_locks_lower_out(51,43);

		normal_cell_50_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,44),
			fetch              => s_fetch(50,44),
			data_in            => s_data_in(50,44),
			data_out           => s_data_out(50,44),
			out1               => s_out1(50,44),
			out2               => s_out2(50,44),
			lock_lower_row_out => s_locks_lower_out(50,44),
			lock_lower_row_in  => s_locks_lower_in(50,44),
			in1                => s_in1(50,44),
			in2                => s_in2(50,44),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(44)
		);
	s_in1(50,44)            <= s_out1(51,44);
	s_in2(50,44)            <= s_out2(51,45);
	s_locks_lower_in(50,44) <= s_locks_lower_out(51,44);

		normal_cell_50_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,45),
			fetch              => s_fetch(50,45),
			data_in            => s_data_in(50,45),
			data_out           => s_data_out(50,45),
			out1               => s_out1(50,45),
			out2               => s_out2(50,45),
			lock_lower_row_out => s_locks_lower_out(50,45),
			lock_lower_row_in  => s_locks_lower_in(50,45),
			in1                => s_in1(50,45),
			in2                => s_in2(50,45),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(45)
		);
	s_in1(50,45)            <= s_out1(51,45);
	s_in2(50,45)            <= s_out2(51,46);
	s_locks_lower_in(50,45) <= s_locks_lower_out(51,45);

		normal_cell_50_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,46),
			fetch              => s_fetch(50,46),
			data_in            => s_data_in(50,46),
			data_out           => s_data_out(50,46),
			out1               => s_out1(50,46),
			out2               => s_out2(50,46),
			lock_lower_row_out => s_locks_lower_out(50,46),
			lock_lower_row_in  => s_locks_lower_in(50,46),
			in1                => s_in1(50,46),
			in2                => s_in2(50,46),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(46)
		);
	s_in1(50,46)            <= s_out1(51,46);
	s_in2(50,46)            <= s_out2(51,47);
	s_locks_lower_in(50,46) <= s_locks_lower_out(51,46);

		normal_cell_50_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,47),
			fetch              => s_fetch(50,47),
			data_in            => s_data_in(50,47),
			data_out           => s_data_out(50,47),
			out1               => s_out1(50,47),
			out2               => s_out2(50,47),
			lock_lower_row_out => s_locks_lower_out(50,47),
			lock_lower_row_in  => s_locks_lower_in(50,47),
			in1                => s_in1(50,47),
			in2                => s_in2(50,47),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(47)
		);
	s_in1(50,47)            <= s_out1(51,47);
	s_in2(50,47)            <= s_out2(51,48);
	s_locks_lower_in(50,47) <= s_locks_lower_out(51,47);

		normal_cell_50_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,48),
			fetch              => s_fetch(50,48),
			data_in            => s_data_in(50,48),
			data_out           => s_data_out(50,48),
			out1               => s_out1(50,48),
			out2               => s_out2(50,48),
			lock_lower_row_out => s_locks_lower_out(50,48),
			lock_lower_row_in  => s_locks_lower_in(50,48),
			in1                => s_in1(50,48),
			in2                => s_in2(50,48),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(48)
		);
	s_in1(50,48)            <= s_out1(51,48);
	s_in2(50,48)            <= s_out2(51,49);
	s_locks_lower_in(50,48) <= s_locks_lower_out(51,48);

		normal_cell_50_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,49),
			fetch              => s_fetch(50,49),
			data_in            => s_data_in(50,49),
			data_out           => s_data_out(50,49),
			out1               => s_out1(50,49),
			out2               => s_out2(50,49),
			lock_lower_row_out => s_locks_lower_out(50,49),
			lock_lower_row_in  => s_locks_lower_in(50,49),
			in1                => s_in1(50,49),
			in2                => s_in2(50,49),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(49)
		);
	s_in1(50,49)            <= s_out1(51,49);
	s_in2(50,49)            <= s_out2(51,50);
	s_locks_lower_in(50,49) <= s_locks_lower_out(51,49);

		normal_cell_50_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,50),
			fetch              => s_fetch(50,50),
			data_in            => s_data_in(50,50),
			data_out           => s_data_out(50,50),
			out1               => s_out1(50,50),
			out2               => s_out2(50,50),
			lock_lower_row_out => s_locks_lower_out(50,50),
			lock_lower_row_in  => s_locks_lower_in(50,50),
			in1                => s_in1(50,50),
			in2                => s_in2(50,50),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(50)
		);
	s_in1(50,50)            <= s_out1(51,50);
	s_in2(50,50)            <= s_out2(51,51);
	s_locks_lower_in(50,50) <= s_locks_lower_out(51,50);

		normal_cell_50_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,51),
			fetch              => s_fetch(50,51),
			data_in            => s_data_in(50,51),
			data_out           => s_data_out(50,51),
			out1               => s_out1(50,51),
			out2               => s_out2(50,51),
			lock_lower_row_out => s_locks_lower_out(50,51),
			lock_lower_row_in  => s_locks_lower_in(50,51),
			in1                => s_in1(50,51),
			in2                => s_in2(50,51),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(51)
		);
	s_in1(50,51)            <= s_out1(51,51);
	s_in2(50,51)            <= s_out2(51,52);
	s_locks_lower_in(50,51) <= s_locks_lower_out(51,51);

		normal_cell_50_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,52),
			fetch              => s_fetch(50,52),
			data_in            => s_data_in(50,52),
			data_out           => s_data_out(50,52),
			out1               => s_out1(50,52),
			out2               => s_out2(50,52),
			lock_lower_row_out => s_locks_lower_out(50,52),
			lock_lower_row_in  => s_locks_lower_in(50,52),
			in1                => s_in1(50,52),
			in2                => s_in2(50,52),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(52)
		);
	s_in1(50,52)            <= s_out1(51,52);
	s_in2(50,52)            <= s_out2(51,53);
	s_locks_lower_in(50,52) <= s_locks_lower_out(51,52);

		normal_cell_50_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,53),
			fetch              => s_fetch(50,53),
			data_in            => s_data_in(50,53),
			data_out           => s_data_out(50,53),
			out1               => s_out1(50,53),
			out2               => s_out2(50,53),
			lock_lower_row_out => s_locks_lower_out(50,53),
			lock_lower_row_in  => s_locks_lower_in(50,53),
			in1                => s_in1(50,53),
			in2                => s_in2(50,53),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(53)
		);
	s_in1(50,53)            <= s_out1(51,53);
	s_in2(50,53)            <= s_out2(51,54);
	s_locks_lower_in(50,53) <= s_locks_lower_out(51,53);

		normal_cell_50_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,54),
			fetch              => s_fetch(50,54),
			data_in            => s_data_in(50,54),
			data_out           => s_data_out(50,54),
			out1               => s_out1(50,54),
			out2               => s_out2(50,54),
			lock_lower_row_out => s_locks_lower_out(50,54),
			lock_lower_row_in  => s_locks_lower_in(50,54),
			in1                => s_in1(50,54),
			in2                => s_in2(50,54),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(54)
		);
	s_in1(50,54)            <= s_out1(51,54);
	s_in2(50,54)            <= s_out2(51,55);
	s_locks_lower_in(50,54) <= s_locks_lower_out(51,54);

		normal_cell_50_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,55),
			fetch              => s_fetch(50,55),
			data_in            => s_data_in(50,55),
			data_out           => s_data_out(50,55),
			out1               => s_out1(50,55),
			out2               => s_out2(50,55),
			lock_lower_row_out => s_locks_lower_out(50,55),
			lock_lower_row_in  => s_locks_lower_in(50,55),
			in1                => s_in1(50,55),
			in2                => s_in2(50,55),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(55)
		);
	s_in1(50,55)            <= s_out1(51,55);
	s_in2(50,55)            <= s_out2(51,56);
	s_locks_lower_in(50,55) <= s_locks_lower_out(51,55);

		normal_cell_50_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,56),
			fetch              => s_fetch(50,56),
			data_in            => s_data_in(50,56),
			data_out           => s_data_out(50,56),
			out1               => s_out1(50,56),
			out2               => s_out2(50,56),
			lock_lower_row_out => s_locks_lower_out(50,56),
			lock_lower_row_in  => s_locks_lower_in(50,56),
			in1                => s_in1(50,56),
			in2                => s_in2(50,56),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(56)
		);
	s_in1(50,56)            <= s_out1(51,56);
	s_in2(50,56)            <= s_out2(51,57);
	s_locks_lower_in(50,56) <= s_locks_lower_out(51,56);

		normal_cell_50_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,57),
			fetch              => s_fetch(50,57),
			data_in            => s_data_in(50,57),
			data_out           => s_data_out(50,57),
			out1               => s_out1(50,57),
			out2               => s_out2(50,57),
			lock_lower_row_out => s_locks_lower_out(50,57),
			lock_lower_row_in  => s_locks_lower_in(50,57),
			in1                => s_in1(50,57),
			in2                => s_in2(50,57),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(57)
		);
	s_in1(50,57)            <= s_out1(51,57);
	s_in2(50,57)            <= s_out2(51,58);
	s_locks_lower_in(50,57) <= s_locks_lower_out(51,57);

		normal_cell_50_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,58),
			fetch              => s_fetch(50,58),
			data_in            => s_data_in(50,58),
			data_out           => s_data_out(50,58),
			out1               => s_out1(50,58),
			out2               => s_out2(50,58),
			lock_lower_row_out => s_locks_lower_out(50,58),
			lock_lower_row_in  => s_locks_lower_in(50,58),
			in1                => s_in1(50,58),
			in2                => s_in2(50,58),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(58)
		);
	s_in1(50,58)            <= s_out1(51,58);
	s_in2(50,58)            <= s_out2(51,59);
	s_locks_lower_in(50,58) <= s_locks_lower_out(51,58);

		normal_cell_50_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,59),
			fetch              => s_fetch(50,59),
			data_in            => s_data_in(50,59),
			data_out           => s_data_out(50,59),
			out1               => s_out1(50,59),
			out2               => s_out2(50,59),
			lock_lower_row_out => s_locks_lower_out(50,59),
			lock_lower_row_in  => s_locks_lower_in(50,59),
			in1                => s_in1(50,59),
			in2                => s_in2(50,59),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(59)
		);
	s_in1(50,59)            <= s_out1(51,59);
	s_in2(50,59)            <= s_out2(51,60);
	s_locks_lower_in(50,59) <= s_locks_lower_out(51,59);

		last_col_cell_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(50,60),
			fetch              => s_fetch(50,60),
			data_in            => s_data_in(50,60),
			data_out           => s_data_out(50,60),
			out1               => s_out1(50,60),
			out2               => s_out2(50,60),
			lock_lower_row_out => s_locks_lower_out(50,60),
			lock_lower_row_in  => s_locks_lower_in(50,60),
			in1                => s_in1(50,60),
			in2                => (others => '0'),
			lock_row           => s_locks(50),
			piv_found          => s_piv_found,
			row_data           => s_row_data(50),
			col_data           => s_col_data(60)
		);
	s_in1(50,60)            <= s_out1(51,60);
	s_locks_lower_in(50,60) <= s_locks_lower_out(51,60);

		normal_cell_51_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,1),
			fetch              => s_fetch(51,1),
			data_in            => s_data_in(51,1),
			data_out           => s_data_out(51,1),
			out1               => s_out1(51,1),
			out2               => s_out2(51,1),
			lock_lower_row_out => s_locks_lower_out(51,1),
			lock_lower_row_in  => s_locks_lower_in(51,1),
			in1                => s_in1(51,1),
			in2                => s_in2(51,1),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(1)
		);
	s_in1(51,1)            <= s_out1(52,1);
	s_in2(51,1)            <= s_out2(52,2);
	s_locks_lower_in(51,1) <= s_locks_lower_out(52,1);

		normal_cell_51_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,2),
			fetch              => s_fetch(51,2),
			data_in            => s_data_in(51,2),
			data_out           => s_data_out(51,2),
			out1               => s_out1(51,2),
			out2               => s_out2(51,2),
			lock_lower_row_out => s_locks_lower_out(51,2),
			lock_lower_row_in  => s_locks_lower_in(51,2),
			in1                => s_in1(51,2),
			in2                => s_in2(51,2),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(2)
		);
	s_in1(51,2)            <= s_out1(52,2);
	s_in2(51,2)            <= s_out2(52,3);
	s_locks_lower_in(51,2) <= s_locks_lower_out(52,2);

		normal_cell_51_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,3),
			fetch              => s_fetch(51,3),
			data_in            => s_data_in(51,3),
			data_out           => s_data_out(51,3),
			out1               => s_out1(51,3),
			out2               => s_out2(51,3),
			lock_lower_row_out => s_locks_lower_out(51,3),
			lock_lower_row_in  => s_locks_lower_in(51,3),
			in1                => s_in1(51,3),
			in2                => s_in2(51,3),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(3)
		);
	s_in1(51,3)            <= s_out1(52,3);
	s_in2(51,3)            <= s_out2(52,4);
	s_locks_lower_in(51,3) <= s_locks_lower_out(52,3);

		normal_cell_51_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,4),
			fetch              => s_fetch(51,4),
			data_in            => s_data_in(51,4),
			data_out           => s_data_out(51,4),
			out1               => s_out1(51,4),
			out2               => s_out2(51,4),
			lock_lower_row_out => s_locks_lower_out(51,4),
			lock_lower_row_in  => s_locks_lower_in(51,4),
			in1                => s_in1(51,4),
			in2                => s_in2(51,4),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(4)
		);
	s_in1(51,4)            <= s_out1(52,4);
	s_in2(51,4)            <= s_out2(52,5);
	s_locks_lower_in(51,4) <= s_locks_lower_out(52,4);

		normal_cell_51_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,5),
			fetch              => s_fetch(51,5),
			data_in            => s_data_in(51,5),
			data_out           => s_data_out(51,5),
			out1               => s_out1(51,5),
			out2               => s_out2(51,5),
			lock_lower_row_out => s_locks_lower_out(51,5),
			lock_lower_row_in  => s_locks_lower_in(51,5),
			in1                => s_in1(51,5),
			in2                => s_in2(51,5),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(5)
		);
	s_in1(51,5)            <= s_out1(52,5);
	s_in2(51,5)            <= s_out2(52,6);
	s_locks_lower_in(51,5) <= s_locks_lower_out(52,5);

		normal_cell_51_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,6),
			fetch              => s_fetch(51,6),
			data_in            => s_data_in(51,6),
			data_out           => s_data_out(51,6),
			out1               => s_out1(51,6),
			out2               => s_out2(51,6),
			lock_lower_row_out => s_locks_lower_out(51,6),
			lock_lower_row_in  => s_locks_lower_in(51,6),
			in1                => s_in1(51,6),
			in2                => s_in2(51,6),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(6)
		);
	s_in1(51,6)            <= s_out1(52,6);
	s_in2(51,6)            <= s_out2(52,7);
	s_locks_lower_in(51,6) <= s_locks_lower_out(52,6);

		normal_cell_51_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,7),
			fetch              => s_fetch(51,7),
			data_in            => s_data_in(51,7),
			data_out           => s_data_out(51,7),
			out1               => s_out1(51,7),
			out2               => s_out2(51,7),
			lock_lower_row_out => s_locks_lower_out(51,7),
			lock_lower_row_in  => s_locks_lower_in(51,7),
			in1                => s_in1(51,7),
			in2                => s_in2(51,7),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(7)
		);
	s_in1(51,7)            <= s_out1(52,7);
	s_in2(51,7)            <= s_out2(52,8);
	s_locks_lower_in(51,7) <= s_locks_lower_out(52,7);

		normal_cell_51_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,8),
			fetch              => s_fetch(51,8),
			data_in            => s_data_in(51,8),
			data_out           => s_data_out(51,8),
			out1               => s_out1(51,8),
			out2               => s_out2(51,8),
			lock_lower_row_out => s_locks_lower_out(51,8),
			lock_lower_row_in  => s_locks_lower_in(51,8),
			in1                => s_in1(51,8),
			in2                => s_in2(51,8),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(8)
		);
	s_in1(51,8)            <= s_out1(52,8);
	s_in2(51,8)            <= s_out2(52,9);
	s_locks_lower_in(51,8) <= s_locks_lower_out(52,8);

		normal_cell_51_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,9),
			fetch              => s_fetch(51,9),
			data_in            => s_data_in(51,9),
			data_out           => s_data_out(51,9),
			out1               => s_out1(51,9),
			out2               => s_out2(51,9),
			lock_lower_row_out => s_locks_lower_out(51,9),
			lock_lower_row_in  => s_locks_lower_in(51,9),
			in1                => s_in1(51,9),
			in2                => s_in2(51,9),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(9)
		);
	s_in1(51,9)            <= s_out1(52,9);
	s_in2(51,9)            <= s_out2(52,10);
	s_locks_lower_in(51,9) <= s_locks_lower_out(52,9);

		normal_cell_51_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,10),
			fetch              => s_fetch(51,10),
			data_in            => s_data_in(51,10),
			data_out           => s_data_out(51,10),
			out1               => s_out1(51,10),
			out2               => s_out2(51,10),
			lock_lower_row_out => s_locks_lower_out(51,10),
			lock_lower_row_in  => s_locks_lower_in(51,10),
			in1                => s_in1(51,10),
			in2                => s_in2(51,10),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(10)
		);
	s_in1(51,10)            <= s_out1(52,10);
	s_in2(51,10)            <= s_out2(52,11);
	s_locks_lower_in(51,10) <= s_locks_lower_out(52,10);

		normal_cell_51_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,11),
			fetch              => s_fetch(51,11),
			data_in            => s_data_in(51,11),
			data_out           => s_data_out(51,11),
			out1               => s_out1(51,11),
			out2               => s_out2(51,11),
			lock_lower_row_out => s_locks_lower_out(51,11),
			lock_lower_row_in  => s_locks_lower_in(51,11),
			in1                => s_in1(51,11),
			in2                => s_in2(51,11),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(11)
		);
	s_in1(51,11)            <= s_out1(52,11);
	s_in2(51,11)            <= s_out2(52,12);
	s_locks_lower_in(51,11) <= s_locks_lower_out(52,11);

		normal_cell_51_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,12),
			fetch              => s_fetch(51,12),
			data_in            => s_data_in(51,12),
			data_out           => s_data_out(51,12),
			out1               => s_out1(51,12),
			out2               => s_out2(51,12),
			lock_lower_row_out => s_locks_lower_out(51,12),
			lock_lower_row_in  => s_locks_lower_in(51,12),
			in1                => s_in1(51,12),
			in2                => s_in2(51,12),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(12)
		);
	s_in1(51,12)            <= s_out1(52,12);
	s_in2(51,12)            <= s_out2(52,13);
	s_locks_lower_in(51,12) <= s_locks_lower_out(52,12);

		normal_cell_51_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,13),
			fetch              => s_fetch(51,13),
			data_in            => s_data_in(51,13),
			data_out           => s_data_out(51,13),
			out1               => s_out1(51,13),
			out2               => s_out2(51,13),
			lock_lower_row_out => s_locks_lower_out(51,13),
			lock_lower_row_in  => s_locks_lower_in(51,13),
			in1                => s_in1(51,13),
			in2                => s_in2(51,13),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(13)
		);
	s_in1(51,13)            <= s_out1(52,13);
	s_in2(51,13)            <= s_out2(52,14);
	s_locks_lower_in(51,13) <= s_locks_lower_out(52,13);

		normal_cell_51_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,14),
			fetch              => s_fetch(51,14),
			data_in            => s_data_in(51,14),
			data_out           => s_data_out(51,14),
			out1               => s_out1(51,14),
			out2               => s_out2(51,14),
			lock_lower_row_out => s_locks_lower_out(51,14),
			lock_lower_row_in  => s_locks_lower_in(51,14),
			in1                => s_in1(51,14),
			in2                => s_in2(51,14),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(14)
		);
	s_in1(51,14)            <= s_out1(52,14);
	s_in2(51,14)            <= s_out2(52,15);
	s_locks_lower_in(51,14) <= s_locks_lower_out(52,14);

		normal_cell_51_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,15),
			fetch              => s_fetch(51,15),
			data_in            => s_data_in(51,15),
			data_out           => s_data_out(51,15),
			out1               => s_out1(51,15),
			out2               => s_out2(51,15),
			lock_lower_row_out => s_locks_lower_out(51,15),
			lock_lower_row_in  => s_locks_lower_in(51,15),
			in1                => s_in1(51,15),
			in2                => s_in2(51,15),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(15)
		);
	s_in1(51,15)            <= s_out1(52,15);
	s_in2(51,15)            <= s_out2(52,16);
	s_locks_lower_in(51,15) <= s_locks_lower_out(52,15);

		normal_cell_51_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,16),
			fetch              => s_fetch(51,16),
			data_in            => s_data_in(51,16),
			data_out           => s_data_out(51,16),
			out1               => s_out1(51,16),
			out2               => s_out2(51,16),
			lock_lower_row_out => s_locks_lower_out(51,16),
			lock_lower_row_in  => s_locks_lower_in(51,16),
			in1                => s_in1(51,16),
			in2                => s_in2(51,16),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(16)
		);
	s_in1(51,16)            <= s_out1(52,16);
	s_in2(51,16)            <= s_out2(52,17);
	s_locks_lower_in(51,16) <= s_locks_lower_out(52,16);

		normal_cell_51_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,17),
			fetch              => s_fetch(51,17),
			data_in            => s_data_in(51,17),
			data_out           => s_data_out(51,17),
			out1               => s_out1(51,17),
			out2               => s_out2(51,17),
			lock_lower_row_out => s_locks_lower_out(51,17),
			lock_lower_row_in  => s_locks_lower_in(51,17),
			in1                => s_in1(51,17),
			in2                => s_in2(51,17),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(17)
		);
	s_in1(51,17)            <= s_out1(52,17);
	s_in2(51,17)            <= s_out2(52,18);
	s_locks_lower_in(51,17) <= s_locks_lower_out(52,17);

		normal_cell_51_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,18),
			fetch              => s_fetch(51,18),
			data_in            => s_data_in(51,18),
			data_out           => s_data_out(51,18),
			out1               => s_out1(51,18),
			out2               => s_out2(51,18),
			lock_lower_row_out => s_locks_lower_out(51,18),
			lock_lower_row_in  => s_locks_lower_in(51,18),
			in1                => s_in1(51,18),
			in2                => s_in2(51,18),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(18)
		);
	s_in1(51,18)            <= s_out1(52,18);
	s_in2(51,18)            <= s_out2(52,19);
	s_locks_lower_in(51,18) <= s_locks_lower_out(52,18);

		normal_cell_51_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,19),
			fetch              => s_fetch(51,19),
			data_in            => s_data_in(51,19),
			data_out           => s_data_out(51,19),
			out1               => s_out1(51,19),
			out2               => s_out2(51,19),
			lock_lower_row_out => s_locks_lower_out(51,19),
			lock_lower_row_in  => s_locks_lower_in(51,19),
			in1                => s_in1(51,19),
			in2                => s_in2(51,19),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(19)
		);
	s_in1(51,19)            <= s_out1(52,19);
	s_in2(51,19)            <= s_out2(52,20);
	s_locks_lower_in(51,19) <= s_locks_lower_out(52,19);

		normal_cell_51_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,20),
			fetch              => s_fetch(51,20),
			data_in            => s_data_in(51,20),
			data_out           => s_data_out(51,20),
			out1               => s_out1(51,20),
			out2               => s_out2(51,20),
			lock_lower_row_out => s_locks_lower_out(51,20),
			lock_lower_row_in  => s_locks_lower_in(51,20),
			in1                => s_in1(51,20),
			in2                => s_in2(51,20),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(20)
		);
	s_in1(51,20)            <= s_out1(52,20);
	s_in2(51,20)            <= s_out2(52,21);
	s_locks_lower_in(51,20) <= s_locks_lower_out(52,20);

		normal_cell_51_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,21),
			fetch              => s_fetch(51,21),
			data_in            => s_data_in(51,21),
			data_out           => s_data_out(51,21),
			out1               => s_out1(51,21),
			out2               => s_out2(51,21),
			lock_lower_row_out => s_locks_lower_out(51,21),
			lock_lower_row_in  => s_locks_lower_in(51,21),
			in1                => s_in1(51,21),
			in2                => s_in2(51,21),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(21)
		);
	s_in1(51,21)            <= s_out1(52,21);
	s_in2(51,21)            <= s_out2(52,22);
	s_locks_lower_in(51,21) <= s_locks_lower_out(52,21);

		normal_cell_51_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,22),
			fetch              => s_fetch(51,22),
			data_in            => s_data_in(51,22),
			data_out           => s_data_out(51,22),
			out1               => s_out1(51,22),
			out2               => s_out2(51,22),
			lock_lower_row_out => s_locks_lower_out(51,22),
			lock_lower_row_in  => s_locks_lower_in(51,22),
			in1                => s_in1(51,22),
			in2                => s_in2(51,22),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(22)
		);
	s_in1(51,22)            <= s_out1(52,22);
	s_in2(51,22)            <= s_out2(52,23);
	s_locks_lower_in(51,22) <= s_locks_lower_out(52,22);

		normal_cell_51_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,23),
			fetch              => s_fetch(51,23),
			data_in            => s_data_in(51,23),
			data_out           => s_data_out(51,23),
			out1               => s_out1(51,23),
			out2               => s_out2(51,23),
			lock_lower_row_out => s_locks_lower_out(51,23),
			lock_lower_row_in  => s_locks_lower_in(51,23),
			in1                => s_in1(51,23),
			in2                => s_in2(51,23),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(23)
		);
	s_in1(51,23)            <= s_out1(52,23);
	s_in2(51,23)            <= s_out2(52,24);
	s_locks_lower_in(51,23) <= s_locks_lower_out(52,23);

		normal_cell_51_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,24),
			fetch              => s_fetch(51,24),
			data_in            => s_data_in(51,24),
			data_out           => s_data_out(51,24),
			out1               => s_out1(51,24),
			out2               => s_out2(51,24),
			lock_lower_row_out => s_locks_lower_out(51,24),
			lock_lower_row_in  => s_locks_lower_in(51,24),
			in1                => s_in1(51,24),
			in2                => s_in2(51,24),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(24)
		);
	s_in1(51,24)            <= s_out1(52,24);
	s_in2(51,24)            <= s_out2(52,25);
	s_locks_lower_in(51,24) <= s_locks_lower_out(52,24);

		normal_cell_51_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,25),
			fetch              => s_fetch(51,25),
			data_in            => s_data_in(51,25),
			data_out           => s_data_out(51,25),
			out1               => s_out1(51,25),
			out2               => s_out2(51,25),
			lock_lower_row_out => s_locks_lower_out(51,25),
			lock_lower_row_in  => s_locks_lower_in(51,25),
			in1                => s_in1(51,25),
			in2                => s_in2(51,25),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(25)
		);
	s_in1(51,25)            <= s_out1(52,25);
	s_in2(51,25)            <= s_out2(52,26);
	s_locks_lower_in(51,25) <= s_locks_lower_out(52,25);

		normal_cell_51_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,26),
			fetch              => s_fetch(51,26),
			data_in            => s_data_in(51,26),
			data_out           => s_data_out(51,26),
			out1               => s_out1(51,26),
			out2               => s_out2(51,26),
			lock_lower_row_out => s_locks_lower_out(51,26),
			lock_lower_row_in  => s_locks_lower_in(51,26),
			in1                => s_in1(51,26),
			in2                => s_in2(51,26),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(26)
		);
	s_in1(51,26)            <= s_out1(52,26);
	s_in2(51,26)            <= s_out2(52,27);
	s_locks_lower_in(51,26) <= s_locks_lower_out(52,26);

		normal_cell_51_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,27),
			fetch              => s_fetch(51,27),
			data_in            => s_data_in(51,27),
			data_out           => s_data_out(51,27),
			out1               => s_out1(51,27),
			out2               => s_out2(51,27),
			lock_lower_row_out => s_locks_lower_out(51,27),
			lock_lower_row_in  => s_locks_lower_in(51,27),
			in1                => s_in1(51,27),
			in2                => s_in2(51,27),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(27)
		);
	s_in1(51,27)            <= s_out1(52,27);
	s_in2(51,27)            <= s_out2(52,28);
	s_locks_lower_in(51,27) <= s_locks_lower_out(52,27);

		normal_cell_51_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,28),
			fetch              => s_fetch(51,28),
			data_in            => s_data_in(51,28),
			data_out           => s_data_out(51,28),
			out1               => s_out1(51,28),
			out2               => s_out2(51,28),
			lock_lower_row_out => s_locks_lower_out(51,28),
			lock_lower_row_in  => s_locks_lower_in(51,28),
			in1                => s_in1(51,28),
			in2                => s_in2(51,28),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(28)
		);
	s_in1(51,28)            <= s_out1(52,28);
	s_in2(51,28)            <= s_out2(52,29);
	s_locks_lower_in(51,28) <= s_locks_lower_out(52,28);

		normal_cell_51_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,29),
			fetch              => s_fetch(51,29),
			data_in            => s_data_in(51,29),
			data_out           => s_data_out(51,29),
			out1               => s_out1(51,29),
			out2               => s_out2(51,29),
			lock_lower_row_out => s_locks_lower_out(51,29),
			lock_lower_row_in  => s_locks_lower_in(51,29),
			in1                => s_in1(51,29),
			in2                => s_in2(51,29),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(29)
		);
	s_in1(51,29)            <= s_out1(52,29);
	s_in2(51,29)            <= s_out2(52,30);
	s_locks_lower_in(51,29) <= s_locks_lower_out(52,29);

		normal_cell_51_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,30),
			fetch              => s_fetch(51,30),
			data_in            => s_data_in(51,30),
			data_out           => s_data_out(51,30),
			out1               => s_out1(51,30),
			out2               => s_out2(51,30),
			lock_lower_row_out => s_locks_lower_out(51,30),
			lock_lower_row_in  => s_locks_lower_in(51,30),
			in1                => s_in1(51,30),
			in2                => s_in2(51,30),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(30)
		);
	s_in1(51,30)            <= s_out1(52,30);
	s_in2(51,30)            <= s_out2(52,31);
	s_locks_lower_in(51,30) <= s_locks_lower_out(52,30);

		normal_cell_51_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,31),
			fetch              => s_fetch(51,31),
			data_in            => s_data_in(51,31),
			data_out           => s_data_out(51,31),
			out1               => s_out1(51,31),
			out2               => s_out2(51,31),
			lock_lower_row_out => s_locks_lower_out(51,31),
			lock_lower_row_in  => s_locks_lower_in(51,31),
			in1                => s_in1(51,31),
			in2                => s_in2(51,31),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(31)
		);
	s_in1(51,31)            <= s_out1(52,31);
	s_in2(51,31)            <= s_out2(52,32);
	s_locks_lower_in(51,31) <= s_locks_lower_out(52,31);

		normal_cell_51_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,32),
			fetch              => s_fetch(51,32),
			data_in            => s_data_in(51,32),
			data_out           => s_data_out(51,32),
			out1               => s_out1(51,32),
			out2               => s_out2(51,32),
			lock_lower_row_out => s_locks_lower_out(51,32),
			lock_lower_row_in  => s_locks_lower_in(51,32),
			in1                => s_in1(51,32),
			in2                => s_in2(51,32),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(32)
		);
	s_in1(51,32)            <= s_out1(52,32);
	s_in2(51,32)            <= s_out2(52,33);
	s_locks_lower_in(51,32) <= s_locks_lower_out(52,32);

		normal_cell_51_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,33),
			fetch              => s_fetch(51,33),
			data_in            => s_data_in(51,33),
			data_out           => s_data_out(51,33),
			out1               => s_out1(51,33),
			out2               => s_out2(51,33),
			lock_lower_row_out => s_locks_lower_out(51,33),
			lock_lower_row_in  => s_locks_lower_in(51,33),
			in1                => s_in1(51,33),
			in2                => s_in2(51,33),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(33)
		);
	s_in1(51,33)            <= s_out1(52,33);
	s_in2(51,33)            <= s_out2(52,34);
	s_locks_lower_in(51,33) <= s_locks_lower_out(52,33);

		normal_cell_51_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,34),
			fetch              => s_fetch(51,34),
			data_in            => s_data_in(51,34),
			data_out           => s_data_out(51,34),
			out1               => s_out1(51,34),
			out2               => s_out2(51,34),
			lock_lower_row_out => s_locks_lower_out(51,34),
			lock_lower_row_in  => s_locks_lower_in(51,34),
			in1                => s_in1(51,34),
			in2                => s_in2(51,34),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(34)
		);
	s_in1(51,34)            <= s_out1(52,34);
	s_in2(51,34)            <= s_out2(52,35);
	s_locks_lower_in(51,34) <= s_locks_lower_out(52,34);

		normal_cell_51_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,35),
			fetch              => s_fetch(51,35),
			data_in            => s_data_in(51,35),
			data_out           => s_data_out(51,35),
			out1               => s_out1(51,35),
			out2               => s_out2(51,35),
			lock_lower_row_out => s_locks_lower_out(51,35),
			lock_lower_row_in  => s_locks_lower_in(51,35),
			in1                => s_in1(51,35),
			in2                => s_in2(51,35),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(35)
		);
	s_in1(51,35)            <= s_out1(52,35);
	s_in2(51,35)            <= s_out2(52,36);
	s_locks_lower_in(51,35) <= s_locks_lower_out(52,35);

		normal_cell_51_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,36),
			fetch              => s_fetch(51,36),
			data_in            => s_data_in(51,36),
			data_out           => s_data_out(51,36),
			out1               => s_out1(51,36),
			out2               => s_out2(51,36),
			lock_lower_row_out => s_locks_lower_out(51,36),
			lock_lower_row_in  => s_locks_lower_in(51,36),
			in1                => s_in1(51,36),
			in2                => s_in2(51,36),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(36)
		);
	s_in1(51,36)            <= s_out1(52,36);
	s_in2(51,36)            <= s_out2(52,37);
	s_locks_lower_in(51,36) <= s_locks_lower_out(52,36);

		normal_cell_51_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,37),
			fetch              => s_fetch(51,37),
			data_in            => s_data_in(51,37),
			data_out           => s_data_out(51,37),
			out1               => s_out1(51,37),
			out2               => s_out2(51,37),
			lock_lower_row_out => s_locks_lower_out(51,37),
			lock_lower_row_in  => s_locks_lower_in(51,37),
			in1                => s_in1(51,37),
			in2                => s_in2(51,37),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(37)
		);
	s_in1(51,37)            <= s_out1(52,37);
	s_in2(51,37)            <= s_out2(52,38);
	s_locks_lower_in(51,37) <= s_locks_lower_out(52,37);

		normal_cell_51_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,38),
			fetch              => s_fetch(51,38),
			data_in            => s_data_in(51,38),
			data_out           => s_data_out(51,38),
			out1               => s_out1(51,38),
			out2               => s_out2(51,38),
			lock_lower_row_out => s_locks_lower_out(51,38),
			lock_lower_row_in  => s_locks_lower_in(51,38),
			in1                => s_in1(51,38),
			in2                => s_in2(51,38),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(38)
		);
	s_in1(51,38)            <= s_out1(52,38);
	s_in2(51,38)            <= s_out2(52,39);
	s_locks_lower_in(51,38) <= s_locks_lower_out(52,38);

		normal_cell_51_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,39),
			fetch              => s_fetch(51,39),
			data_in            => s_data_in(51,39),
			data_out           => s_data_out(51,39),
			out1               => s_out1(51,39),
			out2               => s_out2(51,39),
			lock_lower_row_out => s_locks_lower_out(51,39),
			lock_lower_row_in  => s_locks_lower_in(51,39),
			in1                => s_in1(51,39),
			in2                => s_in2(51,39),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(39)
		);
	s_in1(51,39)            <= s_out1(52,39);
	s_in2(51,39)            <= s_out2(52,40);
	s_locks_lower_in(51,39) <= s_locks_lower_out(52,39);

		normal_cell_51_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,40),
			fetch              => s_fetch(51,40),
			data_in            => s_data_in(51,40),
			data_out           => s_data_out(51,40),
			out1               => s_out1(51,40),
			out2               => s_out2(51,40),
			lock_lower_row_out => s_locks_lower_out(51,40),
			lock_lower_row_in  => s_locks_lower_in(51,40),
			in1                => s_in1(51,40),
			in2                => s_in2(51,40),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(40)
		);
	s_in1(51,40)            <= s_out1(52,40);
	s_in2(51,40)            <= s_out2(52,41);
	s_locks_lower_in(51,40) <= s_locks_lower_out(52,40);

		normal_cell_51_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,41),
			fetch              => s_fetch(51,41),
			data_in            => s_data_in(51,41),
			data_out           => s_data_out(51,41),
			out1               => s_out1(51,41),
			out2               => s_out2(51,41),
			lock_lower_row_out => s_locks_lower_out(51,41),
			lock_lower_row_in  => s_locks_lower_in(51,41),
			in1                => s_in1(51,41),
			in2                => s_in2(51,41),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(41)
		);
	s_in1(51,41)            <= s_out1(52,41);
	s_in2(51,41)            <= s_out2(52,42);
	s_locks_lower_in(51,41) <= s_locks_lower_out(52,41);

		normal_cell_51_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,42),
			fetch              => s_fetch(51,42),
			data_in            => s_data_in(51,42),
			data_out           => s_data_out(51,42),
			out1               => s_out1(51,42),
			out2               => s_out2(51,42),
			lock_lower_row_out => s_locks_lower_out(51,42),
			lock_lower_row_in  => s_locks_lower_in(51,42),
			in1                => s_in1(51,42),
			in2                => s_in2(51,42),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(42)
		);
	s_in1(51,42)            <= s_out1(52,42);
	s_in2(51,42)            <= s_out2(52,43);
	s_locks_lower_in(51,42) <= s_locks_lower_out(52,42);

		normal_cell_51_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,43),
			fetch              => s_fetch(51,43),
			data_in            => s_data_in(51,43),
			data_out           => s_data_out(51,43),
			out1               => s_out1(51,43),
			out2               => s_out2(51,43),
			lock_lower_row_out => s_locks_lower_out(51,43),
			lock_lower_row_in  => s_locks_lower_in(51,43),
			in1                => s_in1(51,43),
			in2                => s_in2(51,43),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(43)
		);
	s_in1(51,43)            <= s_out1(52,43);
	s_in2(51,43)            <= s_out2(52,44);
	s_locks_lower_in(51,43) <= s_locks_lower_out(52,43);

		normal_cell_51_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,44),
			fetch              => s_fetch(51,44),
			data_in            => s_data_in(51,44),
			data_out           => s_data_out(51,44),
			out1               => s_out1(51,44),
			out2               => s_out2(51,44),
			lock_lower_row_out => s_locks_lower_out(51,44),
			lock_lower_row_in  => s_locks_lower_in(51,44),
			in1                => s_in1(51,44),
			in2                => s_in2(51,44),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(44)
		);
	s_in1(51,44)            <= s_out1(52,44);
	s_in2(51,44)            <= s_out2(52,45);
	s_locks_lower_in(51,44) <= s_locks_lower_out(52,44);

		normal_cell_51_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,45),
			fetch              => s_fetch(51,45),
			data_in            => s_data_in(51,45),
			data_out           => s_data_out(51,45),
			out1               => s_out1(51,45),
			out2               => s_out2(51,45),
			lock_lower_row_out => s_locks_lower_out(51,45),
			lock_lower_row_in  => s_locks_lower_in(51,45),
			in1                => s_in1(51,45),
			in2                => s_in2(51,45),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(45)
		);
	s_in1(51,45)            <= s_out1(52,45);
	s_in2(51,45)            <= s_out2(52,46);
	s_locks_lower_in(51,45) <= s_locks_lower_out(52,45);

		normal_cell_51_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,46),
			fetch              => s_fetch(51,46),
			data_in            => s_data_in(51,46),
			data_out           => s_data_out(51,46),
			out1               => s_out1(51,46),
			out2               => s_out2(51,46),
			lock_lower_row_out => s_locks_lower_out(51,46),
			lock_lower_row_in  => s_locks_lower_in(51,46),
			in1                => s_in1(51,46),
			in2                => s_in2(51,46),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(46)
		);
	s_in1(51,46)            <= s_out1(52,46);
	s_in2(51,46)            <= s_out2(52,47);
	s_locks_lower_in(51,46) <= s_locks_lower_out(52,46);

		normal_cell_51_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,47),
			fetch              => s_fetch(51,47),
			data_in            => s_data_in(51,47),
			data_out           => s_data_out(51,47),
			out1               => s_out1(51,47),
			out2               => s_out2(51,47),
			lock_lower_row_out => s_locks_lower_out(51,47),
			lock_lower_row_in  => s_locks_lower_in(51,47),
			in1                => s_in1(51,47),
			in2                => s_in2(51,47),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(47)
		);
	s_in1(51,47)            <= s_out1(52,47);
	s_in2(51,47)            <= s_out2(52,48);
	s_locks_lower_in(51,47) <= s_locks_lower_out(52,47);

		normal_cell_51_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,48),
			fetch              => s_fetch(51,48),
			data_in            => s_data_in(51,48),
			data_out           => s_data_out(51,48),
			out1               => s_out1(51,48),
			out2               => s_out2(51,48),
			lock_lower_row_out => s_locks_lower_out(51,48),
			lock_lower_row_in  => s_locks_lower_in(51,48),
			in1                => s_in1(51,48),
			in2                => s_in2(51,48),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(48)
		);
	s_in1(51,48)            <= s_out1(52,48);
	s_in2(51,48)            <= s_out2(52,49);
	s_locks_lower_in(51,48) <= s_locks_lower_out(52,48);

		normal_cell_51_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,49),
			fetch              => s_fetch(51,49),
			data_in            => s_data_in(51,49),
			data_out           => s_data_out(51,49),
			out1               => s_out1(51,49),
			out2               => s_out2(51,49),
			lock_lower_row_out => s_locks_lower_out(51,49),
			lock_lower_row_in  => s_locks_lower_in(51,49),
			in1                => s_in1(51,49),
			in2                => s_in2(51,49),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(49)
		);
	s_in1(51,49)            <= s_out1(52,49);
	s_in2(51,49)            <= s_out2(52,50);
	s_locks_lower_in(51,49) <= s_locks_lower_out(52,49);

		normal_cell_51_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,50),
			fetch              => s_fetch(51,50),
			data_in            => s_data_in(51,50),
			data_out           => s_data_out(51,50),
			out1               => s_out1(51,50),
			out2               => s_out2(51,50),
			lock_lower_row_out => s_locks_lower_out(51,50),
			lock_lower_row_in  => s_locks_lower_in(51,50),
			in1                => s_in1(51,50),
			in2                => s_in2(51,50),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(50)
		);
	s_in1(51,50)            <= s_out1(52,50);
	s_in2(51,50)            <= s_out2(52,51);
	s_locks_lower_in(51,50) <= s_locks_lower_out(52,50);

		normal_cell_51_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,51),
			fetch              => s_fetch(51,51),
			data_in            => s_data_in(51,51),
			data_out           => s_data_out(51,51),
			out1               => s_out1(51,51),
			out2               => s_out2(51,51),
			lock_lower_row_out => s_locks_lower_out(51,51),
			lock_lower_row_in  => s_locks_lower_in(51,51),
			in1                => s_in1(51,51),
			in2                => s_in2(51,51),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(51)
		);
	s_in1(51,51)            <= s_out1(52,51);
	s_in2(51,51)            <= s_out2(52,52);
	s_locks_lower_in(51,51) <= s_locks_lower_out(52,51);

		normal_cell_51_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,52),
			fetch              => s_fetch(51,52),
			data_in            => s_data_in(51,52),
			data_out           => s_data_out(51,52),
			out1               => s_out1(51,52),
			out2               => s_out2(51,52),
			lock_lower_row_out => s_locks_lower_out(51,52),
			lock_lower_row_in  => s_locks_lower_in(51,52),
			in1                => s_in1(51,52),
			in2                => s_in2(51,52),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(52)
		);
	s_in1(51,52)            <= s_out1(52,52);
	s_in2(51,52)            <= s_out2(52,53);
	s_locks_lower_in(51,52) <= s_locks_lower_out(52,52);

		normal_cell_51_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,53),
			fetch              => s_fetch(51,53),
			data_in            => s_data_in(51,53),
			data_out           => s_data_out(51,53),
			out1               => s_out1(51,53),
			out2               => s_out2(51,53),
			lock_lower_row_out => s_locks_lower_out(51,53),
			lock_lower_row_in  => s_locks_lower_in(51,53),
			in1                => s_in1(51,53),
			in2                => s_in2(51,53),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(53)
		);
	s_in1(51,53)            <= s_out1(52,53);
	s_in2(51,53)            <= s_out2(52,54);
	s_locks_lower_in(51,53) <= s_locks_lower_out(52,53);

		normal_cell_51_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,54),
			fetch              => s_fetch(51,54),
			data_in            => s_data_in(51,54),
			data_out           => s_data_out(51,54),
			out1               => s_out1(51,54),
			out2               => s_out2(51,54),
			lock_lower_row_out => s_locks_lower_out(51,54),
			lock_lower_row_in  => s_locks_lower_in(51,54),
			in1                => s_in1(51,54),
			in2                => s_in2(51,54),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(54)
		);
	s_in1(51,54)            <= s_out1(52,54);
	s_in2(51,54)            <= s_out2(52,55);
	s_locks_lower_in(51,54) <= s_locks_lower_out(52,54);

		normal_cell_51_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,55),
			fetch              => s_fetch(51,55),
			data_in            => s_data_in(51,55),
			data_out           => s_data_out(51,55),
			out1               => s_out1(51,55),
			out2               => s_out2(51,55),
			lock_lower_row_out => s_locks_lower_out(51,55),
			lock_lower_row_in  => s_locks_lower_in(51,55),
			in1                => s_in1(51,55),
			in2                => s_in2(51,55),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(55)
		);
	s_in1(51,55)            <= s_out1(52,55);
	s_in2(51,55)            <= s_out2(52,56);
	s_locks_lower_in(51,55) <= s_locks_lower_out(52,55);

		normal_cell_51_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,56),
			fetch              => s_fetch(51,56),
			data_in            => s_data_in(51,56),
			data_out           => s_data_out(51,56),
			out1               => s_out1(51,56),
			out2               => s_out2(51,56),
			lock_lower_row_out => s_locks_lower_out(51,56),
			lock_lower_row_in  => s_locks_lower_in(51,56),
			in1                => s_in1(51,56),
			in2                => s_in2(51,56),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(56)
		);
	s_in1(51,56)            <= s_out1(52,56);
	s_in2(51,56)            <= s_out2(52,57);
	s_locks_lower_in(51,56) <= s_locks_lower_out(52,56);

		normal_cell_51_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,57),
			fetch              => s_fetch(51,57),
			data_in            => s_data_in(51,57),
			data_out           => s_data_out(51,57),
			out1               => s_out1(51,57),
			out2               => s_out2(51,57),
			lock_lower_row_out => s_locks_lower_out(51,57),
			lock_lower_row_in  => s_locks_lower_in(51,57),
			in1                => s_in1(51,57),
			in2                => s_in2(51,57),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(57)
		);
	s_in1(51,57)            <= s_out1(52,57);
	s_in2(51,57)            <= s_out2(52,58);
	s_locks_lower_in(51,57) <= s_locks_lower_out(52,57);

		normal_cell_51_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,58),
			fetch              => s_fetch(51,58),
			data_in            => s_data_in(51,58),
			data_out           => s_data_out(51,58),
			out1               => s_out1(51,58),
			out2               => s_out2(51,58),
			lock_lower_row_out => s_locks_lower_out(51,58),
			lock_lower_row_in  => s_locks_lower_in(51,58),
			in1                => s_in1(51,58),
			in2                => s_in2(51,58),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(58)
		);
	s_in1(51,58)            <= s_out1(52,58);
	s_in2(51,58)            <= s_out2(52,59);
	s_locks_lower_in(51,58) <= s_locks_lower_out(52,58);

		normal_cell_51_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,59),
			fetch              => s_fetch(51,59),
			data_in            => s_data_in(51,59),
			data_out           => s_data_out(51,59),
			out1               => s_out1(51,59),
			out2               => s_out2(51,59),
			lock_lower_row_out => s_locks_lower_out(51,59),
			lock_lower_row_in  => s_locks_lower_in(51,59),
			in1                => s_in1(51,59),
			in2                => s_in2(51,59),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(59)
		);
	s_in1(51,59)            <= s_out1(52,59);
	s_in2(51,59)            <= s_out2(52,60);
	s_locks_lower_in(51,59) <= s_locks_lower_out(52,59);

		last_col_cell_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(51,60),
			fetch              => s_fetch(51,60),
			data_in            => s_data_in(51,60),
			data_out           => s_data_out(51,60),
			out1               => s_out1(51,60),
			out2               => s_out2(51,60),
			lock_lower_row_out => s_locks_lower_out(51,60),
			lock_lower_row_in  => s_locks_lower_in(51,60),
			in1                => s_in1(51,60),
			in2                => (others => '0'),
			lock_row           => s_locks(51),
			piv_found          => s_piv_found,
			row_data           => s_row_data(51),
			col_data           => s_col_data(60)
		);
	s_in1(51,60)            <= s_out1(52,60);
	s_locks_lower_in(51,60) <= s_locks_lower_out(52,60);

		normal_cell_52_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,1),
			fetch              => s_fetch(52,1),
			data_in            => s_data_in(52,1),
			data_out           => s_data_out(52,1),
			out1               => s_out1(52,1),
			out2               => s_out2(52,1),
			lock_lower_row_out => s_locks_lower_out(52,1),
			lock_lower_row_in  => s_locks_lower_in(52,1),
			in1                => s_in1(52,1),
			in2                => s_in2(52,1),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(1)
		);
	s_in1(52,1)            <= s_out1(53,1);
	s_in2(52,1)            <= s_out2(53,2);
	s_locks_lower_in(52,1) <= s_locks_lower_out(53,1);

		normal_cell_52_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,2),
			fetch              => s_fetch(52,2),
			data_in            => s_data_in(52,2),
			data_out           => s_data_out(52,2),
			out1               => s_out1(52,2),
			out2               => s_out2(52,2),
			lock_lower_row_out => s_locks_lower_out(52,2),
			lock_lower_row_in  => s_locks_lower_in(52,2),
			in1                => s_in1(52,2),
			in2                => s_in2(52,2),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(2)
		);
	s_in1(52,2)            <= s_out1(53,2);
	s_in2(52,2)            <= s_out2(53,3);
	s_locks_lower_in(52,2) <= s_locks_lower_out(53,2);

		normal_cell_52_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,3),
			fetch              => s_fetch(52,3),
			data_in            => s_data_in(52,3),
			data_out           => s_data_out(52,3),
			out1               => s_out1(52,3),
			out2               => s_out2(52,3),
			lock_lower_row_out => s_locks_lower_out(52,3),
			lock_lower_row_in  => s_locks_lower_in(52,3),
			in1                => s_in1(52,3),
			in2                => s_in2(52,3),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(3)
		);
	s_in1(52,3)            <= s_out1(53,3);
	s_in2(52,3)            <= s_out2(53,4);
	s_locks_lower_in(52,3) <= s_locks_lower_out(53,3);

		normal_cell_52_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,4),
			fetch              => s_fetch(52,4),
			data_in            => s_data_in(52,4),
			data_out           => s_data_out(52,4),
			out1               => s_out1(52,4),
			out2               => s_out2(52,4),
			lock_lower_row_out => s_locks_lower_out(52,4),
			lock_lower_row_in  => s_locks_lower_in(52,4),
			in1                => s_in1(52,4),
			in2                => s_in2(52,4),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(4)
		);
	s_in1(52,4)            <= s_out1(53,4);
	s_in2(52,4)            <= s_out2(53,5);
	s_locks_lower_in(52,4) <= s_locks_lower_out(53,4);

		normal_cell_52_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,5),
			fetch              => s_fetch(52,5),
			data_in            => s_data_in(52,5),
			data_out           => s_data_out(52,5),
			out1               => s_out1(52,5),
			out2               => s_out2(52,5),
			lock_lower_row_out => s_locks_lower_out(52,5),
			lock_lower_row_in  => s_locks_lower_in(52,5),
			in1                => s_in1(52,5),
			in2                => s_in2(52,5),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(5)
		);
	s_in1(52,5)            <= s_out1(53,5);
	s_in2(52,5)            <= s_out2(53,6);
	s_locks_lower_in(52,5) <= s_locks_lower_out(53,5);

		normal_cell_52_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,6),
			fetch              => s_fetch(52,6),
			data_in            => s_data_in(52,6),
			data_out           => s_data_out(52,6),
			out1               => s_out1(52,6),
			out2               => s_out2(52,6),
			lock_lower_row_out => s_locks_lower_out(52,6),
			lock_lower_row_in  => s_locks_lower_in(52,6),
			in1                => s_in1(52,6),
			in2                => s_in2(52,6),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(6)
		);
	s_in1(52,6)            <= s_out1(53,6);
	s_in2(52,6)            <= s_out2(53,7);
	s_locks_lower_in(52,6) <= s_locks_lower_out(53,6);

		normal_cell_52_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,7),
			fetch              => s_fetch(52,7),
			data_in            => s_data_in(52,7),
			data_out           => s_data_out(52,7),
			out1               => s_out1(52,7),
			out2               => s_out2(52,7),
			lock_lower_row_out => s_locks_lower_out(52,7),
			lock_lower_row_in  => s_locks_lower_in(52,7),
			in1                => s_in1(52,7),
			in2                => s_in2(52,7),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(7)
		);
	s_in1(52,7)            <= s_out1(53,7);
	s_in2(52,7)            <= s_out2(53,8);
	s_locks_lower_in(52,7) <= s_locks_lower_out(53,7);

		normal_cell_52_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,8),
			fetch              => s_fetch(52,8),
			data_in            => s_data_in(52,8),
			data_out           => s_data_out(52,8),
			out1               => s_out1(52,8),
			out2               => s_out2(52,8),
			lock_lower_row_out => s_locks_lower_out(52,8),
			lock_lower_row_in  => s_locks_lower_in(52,8),
			in1                => s_in1(52,8),
			in2                => s_in2(52,8),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(8)
		);
	s_in1(52,8)            <= s_out1(53,8);
	s_in2(52,8)            <= s_out2(53,9);
	s_locks_lower_in(52,8) <= s_locks_lower_out(53,8);

		normal_cell_52_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,9),
			fetch              => s_fetch(52,9),
			data_in            => s_data_in(52,9),
			data_out           => s_data_out(52,9),
			out1               => s_out1(52,9),
			out2               => s_out2(52,9),
			lock_lower_row_out => s_locks_lower_out(52,9),
			lock_lower_row_in  => s_locks_lower_in(52,9),
			in1                => s_in1(52,9),
			in2                => s_in2(52,9),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(9)
		);
	s_in1(52,9)            <= s_out1(53,9);
	s_in2(52,9)            <= s_out2(53,10);
	s_locks_lower_in(52,9) <= s_locks_lower_out(53,9);

		normal_cell_52_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,10),
			fetch              => s_fetch(52,10),
			data_in            => s_data_in(52,10),
			data_out           => s_data_out(52,10),
			out1               => s_out1(52,10),
			out2               => s_out2(52,10),
			lock_lower_row_out => s_locks_lower_out(52,10),
			lock_lower_row_in  => s_locks_lower_in(52,10),
			in1                => s_in1(52,10),
			in2                => s_in2(52,10),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(10)
		);
	s_in1(52,10)            <= s_out1(53,10);
	s_in2(52,10)            <= s_out2(53,11);
	s_locks_lower_in(52,10) <= s_locks_lower_out(53,10);

		normal_cell_52_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,11),
			fetch              => s_fetch(52,11),
			data_in            => s_data_in(52,11),
			data_out           => s_data_out(52,11),
			out1               => s_out1(52,11),
			out2               => s_out2(52,11),
			lock_lower_row_out => s_locks_lower_out(52,11),
			lock_lower_row_in  => s_locks_lower_in(52,11),
			in1                => s_in1(52,11),
			in2                => s_in2(52,11),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(11)
		);
	s_in1(52,11)            <= s_out1(53,11);
	s_in2(52,11)            <= s_out2(53,12);
	s_locks_lower_in(52,11) <= s_locks_lower_out(53,11);

		normal_cell_52_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,12),
			fetch              => s_fetch(52,12),
			data_in            => s_data_in(52,12),
			data_out           => s_data_out(52,12),
			out1               => s_out1(52,12),
			out2               => s_out2(52,12),
			lock_lower_row_out => s_locks_lower_out(52,12),
			lock_lower_row_in  => s_locks_lower_in(52,12),
			in1                => s_in1(52,12),
			in2                => s_in2(52,12),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(12)
		);
	s_in1(52,12)            <= s_out1(53,12);
	s_in2(52,12)            <= s_out2(53,13);
	s_locks_lower_in(52,12) <= s_locks_lower_out(53,12);

		normal_cell_52_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,13),
			fetch              => s_fetch(52,13),
			data_in            => s_data_in(52,13),
			data_out           => s_data_out(52,13),
			out1               => s_out1(52,13),
			out2               => s_out2(52,13),
			lock_lower_row_out => s_locks_lower_out(52,13),
			lock_lower_row_in  => s_locks_lower_in(52,13),
			in1                => s_in1(52,13),
			in2                => s_in2(52,13),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(13)
		);
	s_in1(52,13)            <= s_out1(53,13);
	s_in2(52,13)            <= s_out2(53,14);
	s_locks_lower_in(52,13) <= s_locks_lower_out(53,13);

		normal_cell_52_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,14),
			fetch              => s_fetch(52,14),
			data_in            => s_data_in(52,14),
			data_out           => s_data_out(52,14),
			out1               => s_out1(52,14),
			out2               => s_out2(52,14),
			lock_lower_row_out => s_locks_lower_out(52,14),
			lock_lower_row_in  => s_locks_lower_in(52,14),
			in1                => s_in1(52,14),
			in2                => s_in2(52,14),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(14)
		);
	s_in1(52,14)            <= s_out1(53,14);
	s_in2(52,14)            <= s_out2(53,15);
	s_locks_lower_in(52,14) <= s_locks_lower_out(53,14);

		normal_cell_52_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,15),
			fetch              => s_fetch(52,15),
			data_in            => s_data_in(52,15),
			data_out           => s_data_out(52,15),
			out1               => s_out1(52,15),
			out2               => s_out2(52,15),
			lock_lower_row_out => s_locks_lower_out(52,15),
			lock_lower_row_in  => s_locks_lower_in(52,15),
			in1                => s_in1(52,15),
			in2                => s_in2(52,15),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(15)
		);
	s_in1(52,15)            <= s_out1(53,15);
	s_in2(52,15)            <= s_out2(53,16);
	s_locks_lower_in(52,15) <= s_locks_lower_out(53,15);

		normal_cell_52_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,16),
			fetch              => s_fetch(52,16),
			data_in            => s_data_in(52,16),
			data_out           => s_data_out(52,16),
			out1               => s_out1(52,16),
			out2               => s_out2(52,16),
			lock_lower_row_out => s_locks_lower_out(52,16),
			lock_lower_row_in  => s_locks_lower_in(52,16),
			in1                => s_in1(52,16),
			in2                => s_in2(52,16),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(16)
		);
	s_in1(52,16)            <= s_out1(53,16);
	s_in2(52,16)            <= s_out2(53,17);
	s_locks_lower_in(52,16) <= s_locks_lower_out(53,16);

		normal_cell_52_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,17),
			fetch              => s_fetch(52,17),
			data_in            => s_data_in(52,17),
			data_out           => s_data_out(52,17),
			out1               => s_out1(52,17),
			out2               => s_out2(52,17),
			lock_lower_row_out => s_locks_lower_out(52,17),
			lock_lower_row_in  => s_locks_lower_in(52,17),
			in1                => s_in1(52,17),
			in2                => s_in2(52,17),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(17)
		);
	s_in1(52,17)            <= s_out1(53,17);
	s_in2(52,17)            <= s_out2(53,18);
	s_locks_lower_in(52,17) <= s_locks_lower_out(53,17);

		normal_cell_52_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,18),
			fetch              => s_fetch(52,18),
			data_in            => s_data_in(52,18),
			data_out           => s_data_out(52,18),
			out1               => s_out1(52,18),
			out2               => s_out2(52,18),
			lock_lower_row_out => s_locks_lower_out(52,18),
			lock_lower_row_in  => s_locks_lower_in(52,18),
			in1                => s_in1(52,18),
			in2                => s_in2(52,18),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(18)
		);
	s_in1(52,18)            <= s_out1(53,18);
	s_in2(52,18)            <= s_out2(53,19);
	s_locks_lower_in(52,18) <= s_locks_lower_out(53,18);

		normal_cell_52_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,19),
			fetch              => s_fetch(52,19),
			data_in            => s_data_in(52,19),
			data_out           => s_data_out(52,19),
			out1               => s_out1(52,19),
			out2               => s_out2(52,19),
			lock_lower_row_out => s_locks_lower_out(52,19),
			lock_lower_row_in  => s_locks_lower_in(52,19),
			in1                => s_in1(52,19),
			in2                => s_in2(52,19),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(19)
		);
	s_in1(52,19)            <= s_out1(53,19);
	s_in2(52,19)            <= s_out2(53,20);
	s_locks_lower_in(52,19) <= s_locks_lower_out(53,19);

		normal_cell_52_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,20),
			fetch              => s_fetch(52,20),
			data_in            => s_data_in(52,20),
			data_out           => s_data_out(52,20),
			out1               => s_out1(52,20),
			out2               => s_out2(52,20),
			lock_lower_row_out => s_locks_lower_out(52,20),
			lock_lower_row_in  => s_locks_lower_in(52,20),
			in1                => s_in1(52,20),
			in2                => s_in2(52,20),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(20)
		);
	s_in1(52,20)            <= s_out1(53,20);
	s_in2(52,20)            <= s_out2(53,21);
	s_locks_lower_in(52,20) <= s_locks_lower_out(53,20);

		normal_cell_52_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,21),
			fetch              => s_fetch(52,21),
			data_in            => s_data_in(52,21),
			data_out           => s_data_out(52,21),
			out1               => s_out1(52,21),
			out2               => s_out2(52,21),
			lock_lower_row_out => s_locks_lower_out(52,21),
			lock_lower_row_in  => s_locks_lower_in(52,21),
			in1                => s_in1(52,21),
			in2                => s_in2(52,21),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(21)
		);
	s_in1(52,21)            <= s_out1(53,21);
	s_in2(52,21)            <= s_out2(53,22);
	s_locks_lower_in(52,21) <= s_locks_lower_out(53,21);

		normal_cell_52_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,22),
			fetch              => s_fetch(52,22),
			data_in            => s_data_in(52,22),
			data_out           => s_data_out(52,22),
			out1               => s_out1(52,22),
			out2               => s_out2(52,22),
			lock_lower_row_out => s_locks_lower_out(52,22),
			lock_lower_row_in  => s_locks_lower_in(52,22),
			in1                => s_in1(52,22),
			in2                => s_in2(52,22),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(22)
		);
	s_in1(52,22)            <= s_out1(53,22);
	s_in2(52,22)            <= s_out2(53,23);
	s_locks_lower_in(52,22) <= s_locks_lower_out(53,22);

		normal_cell_52_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,23),
			fetch              => s_fetch(52,23),
			data_in            => s_data_in(52,23),
			data_out           => s_data_out(52,23),
			out1               => s_out1(52,23),
			out2               => s_out2(52,23),
			lock_lower_row_out => s_locks_lower_out(52,23),
			lock_lower_row_in  => s_locks_lower_in(52,23),
			in1                => s_in1(52,23),
			in2                => s_in2(52,23),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(23)
		);
	s_in1(52,23)            <= s_out1(53,23);
	s_in2(52,23)            <= s_out2(53,24);
	s_locks_lower_in(52,23) <= s_locks_lower_out(53,23);

		normal_cell_52_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,24),
			fetch              => s_fetch(52,24),
			data_in            => s_data_in(52,24),
			data_out           => s_data_out(52,24),
			out1               => s_out1(52,24),
			out2               => s_out2(52,24),
			lock_lower_row_out => s_locks_lower_out(52,24),
			lock_lower_row_in  => s_locks_lower_in(52,24),
			in1                => s_in1(52,24),
			in2                => s_in2(52,24),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(24)
		);
	s_in1(52,24)            <= s_out1(53,24);
	s_in2(52,24)            <= s_out2(53,25);
	s_locks_lower_in(52,24) <= s_locks_lower_out(53,24);

		normal_cell_52_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,25),
			fetch              => s_fetch(52,25),
			data_in            => s_data_in(52,25),
			data_out           => s_data_out(52,25),
			out1               => s_out1(52,25),
			out2               => s_out2(52,25),
			lock_lower_row_out => s_locks_lower_out(52,25),
			lock_lower_row_in  => s_locks_lower_in(52,25),
			in1                => s_in1(52,25),
			in2                => s_in2(52,25),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(25)
		);
	s_in1(52,25)            <= s_out1(53,25);
	s_in2(52,25)            <= s_out2(53,26);
	s_locks_lower_in(52,25) <= s_locks_lower_out(53,25);

		normal_cell_52_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,26),
			fetch              => s_fetch(52,26),
			data_in            => s_data_in(52,26),
			data_out           => s_data_out(52,26),
			out1               => s_out1(52,26),
			out2               => s_out2(52,26),
			lock_lower_row_out => s_locks_lower_out(52,26),
			lock_lower_row_in  => s_locks_lower_in(52,26),
			in1                => s_in1(52,26),
			in2                => s_in2(52,26),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(26)
		);
	s_in1(52,26)            <= s_out1(53,26);
	s_in2(52,26)            <= s_out2(53,27);
	s_locks_lower_in(52,26) <= s_locks_lower_out(53,26);

		normal_cell_52_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,27),
			fetch              => s_fetch(52,27),
			data_in            => s_data_in(52,27),
			data_out           => s_data_out(52,27),
			out1               => s_out1(52,27),
			out2               => s_out2(52,27),
			lock_lower_row_out => s_locks_lower_out(52,27),
			lock_lower_row_in  => s_locks_lower_in(52,27),
			in1                => s_in1(52,27),
			in2                => s_in2(52,27),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(27)
		);
	s_in1(52,27)            <= s_out1(53,27);
	s_in2(52,27)            <= s_out2(53,28);
	s_locks_lower_in(52,27) <= s_locks_lower_out(53,27);

		normal_cell_52_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,28),
			fetch              => s_fetch(52,28),
			data_in            => s_data_in(52,28),
			data_out           => s_data_out(52,28),
			out1               => s_out1(52,28),
			out2               => s_out2(52,28),
			lock_lower_row_out => s_locks_lower_out(52,28),
			lock_lower_row_in  => s_locks_lower_in(52,28),
			in1                => s_in1(52,28),
			in2                => s_in2(52,28),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(28)
		);
	s_in1(52,28)            <= s_out1(53,28);
	s_in2(52,28)            <= s_out2(53,29);
	s_locks_lower_in(52,28) <= s_locks_lower_out(53,28);

		normal_cell_52_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,29),
			fetch              => s_fetch(52,29),
			data_in            => s_data_in(52,29),
			data_out           => s_data_out(52,29),
			out1               => s_out1(52,29),
			out2               => s_out2(52,29),
			lock_lower_row_out => s_locks_lower_out(52,29),
			lock_lower_row_in  => s_locks_lower_in(52,29),
			in1                => s_in1(52,29),
			in2                => s_in2(52,29),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(29)
		);
	s_in1(52,29)            <= s_out1(53,29);
	s_in2(52,29)            <= s_out2(53,30);
	s_locks_lower_in(52,29) <= s_locks_lower_out(53,29);

		normal_cell_52_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,30),
			fetch              => s_fetch(52,30),
			data_in            => s_data_in(52,30),
			data_out           => s_data_out(52,30),
			out1               => s_out1(52,30),
			out2               => s_out2(52,30),
			lock_lower_row_out => s_locks_lower_out(52,30),
			lock_lower_row_in  => s_locks_lower_in(52,30),
			in1                => s_in1(52,30),
			in2                => s_in2(52,30),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(30)
		);
	s_in1(52,30)            <= s_out1(53,30);
	s_in2(52,30)            <= s_out2(53,31);
	s_locks_lower_in(52,30) <= s_locks_lower_out(53,30);

		normal_cell_52_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,31),
			fetch              => s_fetch(52,31),
			data_in            => s_data_in(52,31),
			data_out           => s_data_out(52,31),
			out1               => s_out1(52,31),
			out2               => s_out2(52,31),
			lock_lower_row_out => s_locks_lower_out(52,31),
			lock_lower_row_in  => s_locks_lower_in(52,31),
			in1                => s_in1(52,31),
			in2                => s_in2(52,31),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(31)
		);
	s_in1(52,31)            <= s_out1(53,31);
	s_in2(52,31)            <= s_out2(53,32);
	s_locks_lower_in(52,31) <= s_locks_lower_out(53,31);

		normal_cell_52_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,32),
			fetch              => s_fetch(52,32),
			data_in            => s_data_in(52,32),
			data_out           => s_data_out(52,32),
			out1               => s_out1(52,32),
			out2               => s_out2(52,32),
			lock_lower_row_out => s_locks_lower_out(52,32),
			lock_lower_row_in  => s_locks_lower_in(52,32),
			in1                => s_in1(52,32),
			in2                => s_in2(52,32),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(32)
		);
	s_in1(52,32)            <= s_out1(53,32);
	s_in2(52,32)            <= s_out2(53,33);
	s_locks_lower_in(52,32) <= s_locks_lower_out(53,32);

		normal_cell_52_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,33),
			fetch              => s_fetch(52,33),
			data_in            => s_data_in(52,33),
			data_out           => s_data_out(52,33),
			out1               => s_out1(52,33),
			out2               => s_out2(52,33),
			lock_lower_row_out => s_locks_lower_out(52,33),
			lock_lower_row_in  => s_locks_lower_in(52,33),
			in1                => s_in1(52,33),
			in2                => s_in2(52,33),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(33)
		);
	s_in1(52,33)            <= s_out1(53,33);
	s_in2(52,33)            <= s_out2(53,34);
	s_locks_lower_in(52,33) <= s_locks_lower_out(53,33);

		normal_cell_52_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,34),
			fetch              => s_fetch(52,34),
			data_in            => s_data_in(52,34),
			data_out           => s_data_out(52,34),
			out1               => s_out1(52,34),
			out2               => s_out2(52,34),
			lock_lower_row_out => s_locks_lower_out(52,34),
			lock_lower_row_in  => s_locks_lower_in(52,34),
			in1                => s_in1(52,34),
			in2                => s_in2(52,34),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(34)
		);
	s_in1(52,34)            <= s_out1(53,34);
	s_in2(52,34)            <= s_out2(53,35);
	s_locks_lower_in(52,34) <= s_locks_lower_out(53,34);

		normal_cell_52_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,35),
			fetch              => s_fetch(52,35),
			data_in            => s_data_in(52,35),
			data_out           => s_data_out(52,35),
			out1               => s_out1(52,35),
			out2               => s_out2(52,35),
			lock_lower_row_out => s_locks_lower_out(52,35),
			lock_lower_row_in  => s_locks_lower_in(52,35),
			in1                => s_in1(52,35),
			in2                => s_in2(52,35),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(35)
		);
	s_in1(52,35)            <= s_out1(53,35);
	s_in2(52,35)            <= s_out2(53,36);
	s_locks_lower_in(52,35) <= s_locks_lower_out(53,35);

		normal_cell_52_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,36),
			fetch              => s_fetch(52,36),
			data_in            => s_data_in(52,36),
			data_out           => s_data_out(52,36),
			out1               => s_out1(52,36),
			out2               => s_out2(52,36),
			lock_lower_row_out => s_locks_lower_out(52,36),
			lock_lower_row_in  => s_locks_lower_in(52,36),
			in1                => s_in1(52,36),
			in2                => s_in2(52,36),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(36)
		);
	s_in1(52,36)            <= s_out1(53,36);
	s_in2(52,36)            <= s_out2(53,37);
	s_locks_lower_in(52,36) <= s_locks_lower_out(53,36);

		normal_cell_52_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,37),
			fetch              => s_fetch(52,37),
			data_in            => s_data_in(52,37),
			data_out           => s_data_out(52,37),
			out1               => s_out1(52,37),
			out2               => s_out2(52,37),
			lock_lower_row_out => s_locks_lower_out(52,37),
			lock_lower_row_in  => s_locks_lower_in(52,37),
			in1                => s_in1(52,37),
			in2                => s_in2(52,37),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(37)
		);
	s_in1(52,37)            <= s_out1(53,37);
	s_in2(52,37)            <= s_out2(53,38);
	s_locks_lower_in(52,37) <= s_locks_lower_out(53,37);

		normal_cell_52_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,38),
			fetch              => s_fetch(52,38),
			data_in            => s_data_in(52,38),
			data_out           => s_data_out(52,38),
			out1               => s_out1(52,38),
			out2               => s_out2(52,38),
			lock_lower_row_out => s_locks_lower_out(52,38),
			lock_lower_row_in  => s_locks_lower_in(52,38),
			in1                => s_in1(52,38),
			in2                => s_in2(52,38),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(38)
		);
	s_in1(52,38)            <= s_out1(53,38);
	s_in2(52,38)            <= s_out2(53,39);
	s_locks_lower_in(52,38) <= s_locks_lower_out(53,38);

		normal_cell_52_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,39),
			fetch              => s_fetch(52,39),
			data_in            => s_data_in(52,39),
			data_out           => s_data_out(52,39),
			out1               => s_out1(52,39),
			out2               => s_out2(52,39),
			lock_lower_row_out => s_locks_lower_out(52,39),
			lock_lower_row_in  => s_locks_lower_in(52,39),
			in1                => s_in1(52,39),
			in2                => s_in2(52,39),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(39)
		);
	s_in1(52,39)            <= s_out1(53,39);
	s_in2(52,39)            <= s_out2(53,40);
	s_locks_lower_in(52,39) <= s_locks_lower_out(53,39);

		normal_cell_52_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,40),
			fetch              => s_fetch(52,40),
			data_in            => s_data_in(52,40),
			data_out           => s_data_out(52,40),
			out1               => s_out1(52,40),
			out2               => s_out2(52,40),
			lock_lower_row_out => s_locks_lower_out(52,40),
			lock_lower_row_in  => s_locks_lower_in(52,40),
			in1                => s_in1(52,40),
			in2                => s_in2(52,40),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(40)
		);
	s_in1(52,40)            <= s_out1(53,40);
	s_in2(52,40)            <= s_out2(53,41);
	s_locks_lower_in(52,40) <= s_locks_lower_out(53,40);

		normal_cell_52_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,41),
			fetch              => s_fetch(52,41),
			data_in            => s_data_in(52,41),
			data_out           => s_data_out(52,41),
			out1               => s_out1(52,41),
			out2               => s_out2(52,41),
			lock_lower_row_out => s_locks_lower_out(52,41),
			lock_lower_row_in  => s_locks_lower_in(52,41),
			in1                => s_in1(52,41),
			in2                => s_in2(52,41),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(41)
		);
	s_in1(52,41)            <= s_out1(53,41);
	s_in2(52,41)            <= s_out2(53,42);
	s_locks_lower_in(52,41) <= s_locks_lower_out(53,41);

		normal_cell_52_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,42),
			fetch              => s_fetch(52,42),
			data_in            => s_data_in(52,42),
			data_out           => s_data_out(52,42),
			out1               => s_out1(52,42),
			out2               => s_out2(52,42),
			lock_lower_row_out => s_locks_lower_out(52,42),
			lock_lower_row_in  => s_locks_lower_in(52,42),
			in1                => s_in1(52,42),
			in2                => s_in2(52,42),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(42)
		);
	s_in1(52,42)            <= s_out1(53,42);
	s_in2(52,42)            <= s_out2(53,43);
	s_locks_lower_in(52,42) <= s_locks_lower_out(53,42);

		normal_cell_52_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,43),
			fetch              => s_fetch(52,43),
			data_in            => s_data_in(52,43),
			data_out           => s_data_out(52,43),
			out1               => s_out1(52,43),
			out2               => s_out2(52,43),
			lock_lower_row_out => s_locks_lower_out(52,43),
			lock_lower_row_in  => s_locks_lower_in(52,43),
			in1                => s_in1(52,43),
			in2                => s_in2(52,43),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(43)
		);
	s_in1(52,43)            <= s_out1(53,43);
	s_in2(52,43)            <= s_out2(53,44);
	s_locks_lower_in(52,43) <= s_locks_lower_out(53,43);

		normal_cell_52_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,44),
			fetch              => s_fetch(52,44),
			data_in            => s_data_in(52,44),
			data_out           => s_data_out(52,44),
			out1               => s_out1(52,44),
			out2               => s_out2(52,44),
			lock_lower_row_out => s_locks_lower_out(52,44),
			lock_lower_row_in  => s_locks_lower_in(52,44),
			in1                => s_in1(52,44),
			in2                => s_in2(52,44),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(44)
		);
	s_in1(52,44)            <= s_out1(53,44);
	s_in2(52,44)            <= s_out2(53,45);
	s_locks_lower_in(52,44) <= s_locks_lower_out(53,44);

		normal_cell_52_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,45),
			fetch              => s_fetch(52,45),
			data_in            => s_data_in(52,45),
			data_out           => s_data_out(52,45),
			out1               => s_out1(52,45),
			out2               => s_out2(52,45),
			lock_lower_row_out => s_locks_lower_out(52,45),
			lock_lower_row_in  => s_locks_lower_in(52,45),
			in1                => s_in1(52,45),
			in2                => s_in2(52,45),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(45)
		);
	s_in1(52,45)            <= s_out1(53,45);
	s_in2(52,45)            <= s_out2(53,46);
	s_locks_lower_in(52,45) <= s_locks_lower_out(53,45);

		normal_cell_52_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,46),
			fetch              => s_fetch(52,46),
			data_in            => s_data_in(52,46),
			data_out           => s_data_out(52,46),
			out1               => s_out1(52,46),
			out2               => s_out2(52,46),
			lock_lower_row_out => s_locks_lower_out(52,46),
			lock_lower_row_in  => s_locks_lower_in(52,46),
			in1                => s_in1(52,46),
			in2                => s_in2(52,46),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(46)
		);
	s_in1(52,46)            <= s_out1(53,46);
	s_in2(52,46)            <= s_out2(53,47);
	s_locks_lower_in(52,46) <= s_locks_lower_out(53,46);

		normal_cell_52_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,47),
			fetch              => s_fetch(52,47),
			data_in            => s_data_in(52,47),
			data_out           => s_data_out(52,47),
			out1               => s_out1(52,47),
			out2               => s_out2(52,47),
			lock_lower_row_out => s_locks_lower_out(52,47),
			lock_lower_row_in  => s_locks_lower_in(52,47),
			in1                => s_in1(52,47),
			in2                => s_in2(52,47),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(47)
		);
	s_in1(52,47)            <= s_out1(53,47);
	s_in2(52,47)            <= s_out2(53,48);
	s_locks_lower_in(52,47) <= s_locks_lower_out(53,47);

		normal_cell_52_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,48),
			fetch              => s_fetch(52,48),
			data_in            => s_data_in(52,48),
			data_out           => s_data_out(52,48),
			out1               => s_out1(52,48),
			out2               => s_out2(52,48),
			lock_lower_row_out => s_locks_lower_out(52,48),
			lock_lower_row_in  => s_locks_lower_in(52,48),
			in1                => s_in1(52,48),
			in2                => s_in2(52,48),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(48)
		);
	s_in1(52,48)            <= s_out1(53,48);
	s_in2(52,48)            <= s_out2(53,49);
	s_locks_lower_in(52,48) <= s_locks_lower_out(53,48);

		normal_cell_52_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,49),
			fetch              => s_fetch(52,49),
			data_in            => s_data_in(52,49),
			data_out           => s_data_out(52,49),
			out1               => s_out1(52,49),
			out2               => s_out2(52,49),
			lock_lower_row_out => s_locks_lower_out(52,49),
			lock_lower_row_in  => s_locks_lower_in(52,49),
			in1                => s_in1(52,49),
			in2                => s_in2(52,49),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(49)
		);
	s_in1(52,49)            <= s_out1(53,49);
	s_in2(52,49)            <= s_out2(53,50);
	s_locks_lower_in(52,49) <= s_locks_lower_out(53,49);

		normal_cell_52_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,50),
			fetch              => s_fetch(52,50),
			data_in            => s_data_in(52,50),
			data_out           => s_data_out(52,50),
			out1               => s_out1(52,50),
			out2               => s_out2(52,50),
			lock_lower_row_out => s_locks_lower_out(52,50),
			lock_lower_row_in  => s_locks_lower_in(52,50),
			in1                => s_in1(52,50),
			in2                => s_in2(52,50),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(50)
		);
	s_in1(52,50)            <= s_out1(53,50);
	s_in2(52,50)            <= s_out2(53,51);
	s_locks_lower_in(52,50) <= s_locks_lower_out(53,50);

		normal_cell_52_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,51),
			fetch              => s_fetch(52,51),
			data_in            => s_data_in(52,51),
			data_out           => s_data_out(52,51),
			out1               => s_out1(52,51),
			out2               => s_out2(52,51),
			lock_lower_row_out => s_locks_lower_out(52,51),
			lock_lower_row_in  => s_locks_lower_in(52,51),
			in1                => s_in1(52,51),
			in2                => s_in2(52,51),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(51)
		);
	s_in1(52,51)            <= s_out1(53,51);
	s_in2(52,51)            <= s_out2(53,52);
	s_locks_lower_in(52,51) <= s_locks_lower_out(53,51);

		normal_cell_52_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,52),
			fetch              => s_fetch(52,52),
			data_in            => s_data_in(52,52),
			data_out           => s_data_out(52,52),
			out1               => s_out1(52,52),
			out2               => s_out2(52,52),
			lock_lower_row_out => s_locks_lower_out(52,52),
			lock_lower_row_in  => s_locks_lower_in(52,52),
			in1                => s_in1(52,52),
			in2                => s_in2(52,52),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(52)
		);
	s_in1(52,52)            <= s_out1(53,52);
	s_in2(52,52)            <= s_out2(53,53);
	s_locks_lower_in(52,52) <= s_locks_lower_out(53,52);

		normal_cell_52_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,53),
			fetch              => s_fetch(52,53),
			data_in            => s_data_in(52,53),
			data_out           => s_data_out(52,53),
			out1               => s_out1(52,53),
			out2               => s_out2(52,53),
			lock_lower_row_out => s_locks_lower_out(52,53),
			lock_lower_row_in  => s_locks_lower_in(52,53),
			in1                => s_in1(52,53),
			in2                => s_in2(52,53),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(53)
		);
	s_in1(52,53)            <= s_out1(53,53);
	s_in2(52,53)            <= s_out2(53,54);
	s_locks_lower_in(52,53) <= s_locks_lower_out(53,53);

		normal_cell_52_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,54),
			fetch              => s_fetch(52,54),
			data_in            => s_data_in(52,54),
			data_out           => s_data_out(52,54),
			out1               => s_out1(52,54),
			out2               => s_out2(52,54),
			lock_lower_row_out => s_locks_lower_out(52,54),
			lock_lower_row_in  => s_locks_lower_in(52,54),
			in1                => s_in1(52,54),
			in2                => s_in2(52,54),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(54)
		);
	s_in1(52,54)            <= s_out1(53,54);
	s_in2(52,54)            <= s_out2(53,55);
	s_locks_lower_in(52,54) <= s_locks_lower_out(53,54);

		normal_cell_52_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,55),
			fetch              => s_fetch(52,55),
			data_in            => s_data_in(52,55),
			data_out           => s_data_out(52,55),
			out1               => s_out1(52,55),
			out2               => s_out2(52,55),
			lock_lower_row_out => s_locks_lower_out(52,55),
			lock_lower_row_in  => s_locks_lower_in(52,55),
			in1                => s_in1(52,55),
			in2                => s_in2(52,55),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(55)
		);
	s_in1(52,55)            <= s_out1(53,55);
	s_in2(52,55)            <= s_out2(53,56);
	s_locks_lower_in(52,55) <= s_locks_lower_out(53,55);

		normal_cell_52_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,56),
			fetch              => s_fetch(52,56),
			data_in            => s_data_in(52,56),
			data_out           => s_data_out(52,56),
			out1               => s_out1(52,56),
			out2               => s_out2(52,56),
			lock_lower_row_out => s_locks_lower_out(52,56),
			lock_lower_row_in  => s_locks_lower_in(52,56),
			in1                => s_in1(52,56),
			in2                => s_in2(52,56),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(56)
		);
	s_in1(52,56)            <= s_out1(53,56);
	s_in2(52,56)            <= s_out2(53,57);
	s_locks_lower_in(52,56) <= s_locks_lower_out(53,56);

		normal_cell_52_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,57),
			fetch              => s_fetch(52,57),
			data_in            => s_data_in(52,57),
			data_out           => s_data_out(52,57),
			out1               => s_out1(52,57),
			out2               => s_out2(52,57),
			lock_lower_row_out => s_locks_lower_out(52,57),
			lock_lower_row_in  => s_locks_lower_in(52,57),
			in1                => s_in1(52,57),
			in2                => s_in2(52,57),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(57)
		);
	s_in1(52,57)            <= s_out1(53,57);
	s_in2(52,57)            <= s_out2(53,58);
	s_locks_lower_in(52,57) <= s_locks_lower_out(53,57);

		normal_cell_52_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,58),
			fetch              => s_fetch(52,58),
			data_in            => s_data_in(52,58),
			data_out           => s_data_out(52,58),
			out1               => s_out1(52,58),
			out2               => s_out2(52,58),
			lock_lower_row_out => s_locks_lower_out(52,58),
			lock_lower_row_in  => s_locks_lower_in(52,58),
			in1                => s_in1(52,58),
			in2                => s_in2(52,58),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(58)
		);
	s_in1(52,58)            <= s_out1(53,58);
	s_in2(52,58)            <= s_out2(53,59);
	s_locks_lower_in(52,58) <= s_locks_lower_out(53,58);

		normal_cell_52_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,59),
			fetch              => s_fetch(52,59),
			data_in            => s_data_in(52,59),
			data_out           => s_data_out(52,59),
			out1               => s_out1(52,59),
			out2               => s_out2(52,59),
			lock_lower_row_out => s_locks_lower_out(52,59),
			lock_lower_row_in  => s_locks_lower_in(52,59),
			in1                => s_in1(52,59),
			in2                => s_in2(52,59),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(59)
		);
	s_in1(52,59)            <= s_out1(53,59);
	s_in2(52,59)            <= s_out2(53,60);
	s_locks_lower_in(52,59) <= s_locks_lower_out(53,59);

		last_col_cell_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(52,60),
			fetch              => s_fetch(52,60),
			data_in            => s_data_in(52,60),
			data_out           => s_data_out(52,60),
			out1               => s_out1(52,60),
			out2               => s_out2(52,60),
			lock_lower_row_out => s_locks_lower_out(52,60),
			lock_lower_row_in  => s_locks_lower_in(52,60),
			in1                => s_in1(52,60),
			in2                => (others => '0'),
			lock_row           => s_locks(52),
			piv_found          => s_piv_found,
			row_data           => s_row_data(52),
			col_data           => s_col_data(60)
		);
	s_in1(52,60)            <= s_out1(53,60);
	s_locks_lower_in(52,60) <= s_locks_lower_out(53,60);

		normal_cell_53_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,1),
			fetch              => s_fetch(53,1),
			data_in            => s_data_in(53,1),
			data_out           => s_data_out(53,1),
			out1               => s_out1(53,1),
			out2               => s_out2(53,1),
			lock_lower_row_out => s_locks_lower_out(53,1),
			lock_lower_row_in  => s_locks_lower_in(53,1),
			in1                => s_in1(53,1),
			in2                => s_in2(53,1),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(1)
		);
	s_in1(53,1)            <= s_out1(54,1);
	s_in2(53,1)            <= s_out2(54,2);
	s_locks_lower_in(53,1) <= s_locks_lower_out(54,1);

		normal_cell_53_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,2),
			fetch              => s_fetch(53,2),
			data_in            => s_data_in(53,2),
			data_out           => s_data_out(53,2),
			out1               => s_out1(53,2),
			out2               => s_out2(53,2),
			lock_lower_row_out => s_locks_lower_out(53,2),
			lock_lower_row_in  => s_locks_lower_in(53,2),
			in1                => s_in1(53,2),
			in2                => s_in2(53,2),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(2)
		);
	s_in1(53,2)            <= s_out1(54,2);
	s_in2(53,2)            <= s_out2(54,3);
	s_locks_lower_in(53,2) <= s_locks_lower_out(54,2);

		normal_cell_53_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,3),
			fetch              => s_fetch(53,3),
			data_in            => s_data_in(53,3),
			data_out           => s_data_out(53,3),
			out1               => s_out1(53,3),
			out2               => s_out2(53,3),
			lock_lower_row_out => s_locks_lower_out(53,3),
			lock_lower_row_in  => s_locks_lower_in(53,3),
			in1                => s_in1(53,3),
			in2                => s_in2(53,3),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(3)
		);
	s_in1(53,3)            <= s_out1(54,3);
	s_in2(53,3)            <= s_out2(54,4);
	s_locks_lower_in(53,3) <= s_locks_lower_out(54,3);

		normal_cell_53_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,4),
			fetch              => s_fetch(53,4),
			data_in            => s_data_in(53,4),
			data_out           => s_data_out(53,4),
			out1               => s_out1(53,4),
			out2               => s_out2(53,4),
			lock_lower_row_out => s_locks_lower_out(53,4),
			lock_lower_row_in  => s_locks_lower_in(53,4),
			in1                => s_in1(53,4),
			in2                => s_in2(53,4),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(4)
		);
	s_in1(53,4)            <= s_out1(54,4);
	s_in2(53,4)            <= s_out2(54,5);
	s_locks_lower_in(53,4) <= s_locks_lower_out(54,4);

		normal_cell_53_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,5),
			fetch              => s_fetch(53,5),
			data_in            => s_data_in(53,5),
			data_out           => s_data_out(53,5),
			out1               => s_out1(53,5),
			out2               => s_out2(53,5),
			lock_lower_row_out => s_locks_lower_out(53,5),
			lock_lower_row_in  => s_locks_lower_in(53,5),
			in1                => s_in1(53,5),
			in2                => s_in2(53,5),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(5)
		);
	s_in1(53,5)            <= s_out1(54,5);
	s_in2(53,5)            <= s_out2(54,6);
	s_locks_lower_in(53,5) <= s_locks_lower_out(54,5);

		normal_cell_53_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,6),
			fetch              => s_fetch(53,6),
			data_in            => s_data_in(53,6),
			data_out           => s_data_out(53,6),
			out1               => s_out1(53,6),
			out2               => s_out2(53,6),
			lock_lower_row_out => s_locks_lower_out(53,6),
			lock_lower_row_in  => s_locks_lower_in(53,6),
			in1                => s_in1(53,6),
			in2                => s_in2(53,6),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(6)
		);
	s_in1(53,6)            <= s_out1(54,6);
	s_in2(53,6)            <= s_out2(54,7);
	s_locks_lower_in(53,6) <= s_locks_lower_out(54,6);

		normal_cell_53_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,7),
			fetch              => s_fetch(53,7),
			data_in            => s_data_in(53,7),
			data_out           => s_data_out(53,7),
			out1               => s_out1(53,7),
			out2               => s_out2(53,7),
			lock_lower_row_out => s_locks_lower_out(53,7),
			lock_lower_row_in  => s_locks_lower_in(53,7),
			in1                => s_in1(53,7),
			in2                => s_in2(53,7),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(7)
		);
	s_in1(53,7)            <= s_out1(54,7);
	s_in2(53,7)            <= s_out2(54,8);
	s_locks_lower_in(53,7) <= s_locks_lower_out(54,7);

		normal_cell_53_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,8),
			fetch              => s_fetch(53,8),
			data_in            => s_data_in(53,8),
			data_out           => s_data_out(53,8),
			out1               => s_out1(53,8),
			out2               => s_out2(53,8),
			lock_lower_row_out => s_locks_lower_out(53,8),
			lock_lower_row_in  => s_locks_lower_in(53,8),
			in1                => s_in1(53,8),
			in2                => s_in2(53,8),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(8)
		);
	s_in1(53,8)            <= s_out1(54,8);
	s_in2(53,8)            <= s_out2(54,9);
	s_locks_lower_in(53,8) <= s_locks_lower_out(54,8);

		normal_cell_53_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,9),
			fetch              => s_fetch(53,9),
			data_in            => s_data_in(53,9),
			data_out           => s_data_out(53,9),
			out1               => s_out1(53,9),
			out2               => s_out2(53,9),
			lock_lower_row_out => s_locks_lower_out(53,9),
			lock_lower_row_in  => s_locks_lower_in(53,9),
			in1                => s_in1(53,9),
			in2                => s_in2(53,9),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(9)
		);
	s_in1(53,9)            <= s_out1(54,9);
	s_in2(53,9)            <= s_out2(54,10);
	s_locks_lower_in(53,9) <= s_locks_lower_out(54,9);

		normal_cell_53_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,10),
			fetch              => s_fetch(53,10),
			data_in            => s_data_in(53,10),
			data_out           => s_data_out(53,10),
			out1               => s_out1(53,10),
			out2               => s_out2(53,10),
			lock_lower_row_out => s_locks_lower_out(53,10),
			lock_lower_row_in  => s_locks_lower_in(53,10),
			in1                => s_in1(53,10),
			in2                => s_in2(53,10),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(10)
		);
	s_in1(53,10)            <= s_out1(54,10);
	s_in2(53,10)            <= s_out2(54,11);
	s_locks_lower_in(53,10) <= s_locks_lower_out(54,10);

		normal_cell_53_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,11),
			fetch              => s_fetch(53,11),
			data_in            => s_data_in(53,11),
			data_out           => s_data_out(53,11),
			out1               => s_out1(53,11),
			out2               => s_out2(53,11),
			lock_lower_row_out => s_locks_lower_out(53,11),
			lock_lower_row_in  => s_locks_lower_in(53,11),
			in1                => s_in1(53,11),
			in2                => s_in2(53,11),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(11)
		);
	s_in1(53,11)            <= s_out1(54,11);
	s_in2(53,11)            <= s_out2(54,12);
	s_locks_lower_in(53,11) <= s_locks_lower_out(54,11);

		normal_cell_53_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,12),
			fetch              => s_fetch(53,12),
			data_in            => s_data_in(53,12),
			data_out           => s_data_out(53,12),
			out1               => s_out1(53,12),
			out2               => s_out2(53,12),
			lock_lower_row_out => s_locks_lower_out(53,12),
			lock_lower_row_in  => s_locks_lower_in(53,12),
			in1                => s_in1(53,12),
			in2                => s_in2(53,12),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(12)
		);
	s_in1(53,12)            <= s_out1(54,12);
	s_in2(53,12)            <= s_out2(54,13);
	s_locks_lower_in(53,12) <= s_locks_lower_out(54,12);

		normal_cell_53_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,13),
			fetch              => s_fetch(53,13),
			data_in            => s_data_in(53,13),
			data_out           => s_data_out(53,13),
			out1               => s_out1(53,13),
			out2               => s_out2(53,13),
			lock_lower_row_out => s_locks_lower_out(53,13),
			lock_lower_row_in  => s_locks_lower_in(53,13),
			in1                => s_in1(53,13),
			in2                => s_in2(53,13),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(13)
		);
	s_in1(53,13)            <= s_out1(54,13);
	s_in2(53,13)            <= s_out2(54,14);
	s_locks_lower_in(53,13) <= s_locks_lower_out(54,13);

		normal_cell_53_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,14),
			fetch              => s_fetch(53,14),
			data_in            => s_data_in(53,14),
			data_out           => s_data_out(53,14),
			out1               => s_out1(53,14),
			out2               => s_out2(53,14),
			lock_lower_row_out => s_locks_lower_out(53,14),
			lock_lower_row_in  => s_locks_lower_in(53,14),
			in1                => s_in1(53,14),
			in2                => s_in2(53,14),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(14)
		);
	s_in1(53,14)            <= s_out1(54,14);
	s_in2(53,14)            <= s_out2(54,15);
	s_locks_lower_in(53,14) <= s_locks_lower_out(54,14);

		normal_cell_53_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,15),
			fetch              => s_fetch(53,15),
			data_in            => s_data_in(53,15),
			data_out           => s_data_out(53,15),
			out1               => s_out1(53,15),
			out2               => s_out2(53,15),
			lock_lower_row_out => s_locks_lower_out(53,15),
			lock_lower_row_in  => s_locks_lower_in(53,15),
			in1                => s_in1(53,15),
			in2                => s_in2(53,15),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(15)
		);
	s_in1(53,15)            <= s_out1(54,15);
	s_in2(53,15)            <= s_out2(54,16);
	s_locks_lower_in(53,15) <= s_locks_lower_out(54,15);

		normal_cell_53_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,16),
			fetch              => s_fetch(53,16),
			data_in            => s_data_in(53,16),
			data_out           => s_data_out(53,16),
			out1               => s_out1(53,16),
			out2               => s_out2(53,16),
			lock_lower_row_out => s_locks_lower_out(53,16),
			lock_lower_row_in  => s_locks_lower_in(53,16),
			in1                => s_in1(53,16),
			in2                => s_in2(53,16),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(16)
		);
	s_in1(53,16)            <= s_out1(54,16);
	s_in2(53,16)            <= s_out2(54,17);
	s_locks_lower_in(53,16) <= s_locks_lower_out(54,16);

		normal_cell_53_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,17),
			fetch              => s_fetch(53,17),
			data_in            => s_data_in(53,17),
			data_out           => s_data_out(53,17),
			out1               => s_out1(53,17),
			out2               => s_out2(53,17),
			lock_lower_row_out => s_locks_lower_out(53,17),
			lock_lower_row_in  => s_locks_lower_in(53,17),
			in1                => s_in1(53,17),
			in2                => s_in2(53,17),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(17)
		);
	s_in1(53,17)            <= s_out1(54,17);
	s_in2(53,17)            <= s_out2(54,18);
	s_locks_lower_in(53,17) <= s_locks_lower_out(54,17);

		normal_cell_53_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,18),
			fetch              => s_fetch(53,18),
			data_in            => s_data_in(53,18),
			data_out           => s_data_out(53,18),
			out1               => s_out1(53,18),
			out2               => s_out2(53,18),
			lock_lower_row_out => s_locks_lower_out(53,18),
			lock_lower_row_in  => s_locks_lower_in(53,18),
			in1                => s_in1(53,18),
			in2                => s_in2(53,18),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(18)
		);
	s_in1(53,18)            <= s_out1(54,18);
	s_in2(53,18)            <= s_out2(54,19);
	s_locks_lower_in(53,18) <= s_locks_lower_out(54,18);

		normal_cell_53_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,19),
			fetch              => s_fetch(53,19),
			data_in            => s_data_in(53,19),
			data_out           => s_data_out(53,19),
			out1               => s_out1(53,19),
			out2               => s_out2(53,19),
			lock_lower_row_out => s_locks_lower_out(53,19),
			lock_lower_row_in  => s_locks_lower_in(53,19),
			in1                => s_in1(53,19),
			in2                => s_in2(53,19),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(19)
		);
	s_in1(53,19)            <= s_out1(54,19);
	s_in2(53,19)            <= s_out2(54,20);
	s_locks_lower_in(53,19) <= s_locks_lower_out(54,19);

		normal_cell_53_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,20),
			fetch              => s_fetch(53,20),
			data_in            => s_data_in(53,20),
			data_out           => s_data_out(53,20),
			out1               => s_out1(53,20),
			out2               => s_out2(53,20),
			lock_lower_row_out => s_locks_lower_out(53,20),
			lock_lower_row_in  => s_locks_lower_in(53,20),
			in1                => s_in1(53,20),
			in2                => s_in2(53,20),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(20)
		);
	s_in1(53,20)            <= s_out1(54,20);
	s_in2(53,20)            <= s_out2(54,21);
	s_locks_lower_in(53,20) <= s_locks_lower_out(54,20);

		normal_cell_53_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,21),
			fetch              => s_fetch(53,21),
			data_in            => s_data_in(53,21),
			data_out           => s_data_out(53,21),
			out1               => s_out1(53,21),
			out2               => s_out2(53,21),
			lock_lower_row_out => s_locks_lower_out(53,21),
			lock_lower_row_in  => s_locks_lower_in(53,21),
			in1                => s_in1(53,21),
			in2                => s_in2(53,21),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(21)
		);
	s_in1(53,21)            <= s_out1(54,21);
	s_in2(53,21)            <= s_out2(54,22);
	s_locks_lower_in(53,21) <= s_locks_lower_out(54,21);

		normal_cell_53_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,22),
			fetch              => s_fetch(53,22),
			data_in            => s_data_in(53,22),
			data_out           => s_data_out(53,22),
			out1               => s_out1(53,22),
			out2               => s_out2(53,22),
			lock_lower_row_out => s_locks_lower_out(53,22),
			lock_lower_row_in  => s_locks_lower_in(53,22),
			in1                => s_in1(53,22),
			in2                => s_in2(53,22),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(22)
		);
	s_in1(53,22)            <= s_out1(54,22);
	s_in2(53,22)            <= s_out2(54,23);
	s_locks_lower_in(53,22) <= s_locks_lower_out(54,22);

		normal_cell_53_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,23),
			fetch              => s_fetch(53,23),
			data_in            => s_data_in(53,23),
			data_out           => s_data_out(53,23),
			out1               => s_out1(53,23),
			out2               => s_out2(53,23),
			lock_lower_row_out => s_locks_lower_out(53,23),
			lock_lower_row_in  => s_locks_lower_in(53,23),
			in1                => s_in1(53,23),
			in2                => s_in2(53,23),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(23)
		);
	s_in1(53,23)            <= s_out1(54,23);
	s_in2(53,23)            <= s_out2(54,24);
	s_locks_lower_in(53,23) <= s_locks_lower_out(54,23);

		normal_cell_53_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,24),
			fetch              => s_fetch(53,24),
			data_in            => s_data_in(53,24),
			data_out           => s_data_out(53,24),
			out1               => s_out1(53,24),
			out2               => s_out2(53,24),
			lock_lower_row_out => s_locks_lower_out(53,24),
			lock_lower_row_in  => s_locks_lower_in(53,24),
			in1                => s_in1(53,24),
			in2                => s_in2(53,24),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(24)
		);
	s_in1(53,24)            <= s_out1(54,24);
	s_in2(53,24)            <= s_out2(54,25);
	s_locks_lower_in(53,24) <= s_locks_lower_out(54,24);

		normal_cell_53_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,25),
			fetch              => s_fetch(53,25),
			data_in            => s_data_in(53,25),
			data_out           => s_data_out(53,25),
			out1               => s_out1(53,25),
			out2               => s_out2(53,25),
			lock_lower_row_out => s_locks_lower_out(53,25),
			lock_lower_row_in  => s_locks_lower_in(53,25),
			in1                => s_in1(53,25),
			in2                => s_in2(53,25),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(25)
		);
	s_in1(53,25)            <= s_out1(54,25);
	s_in2(53,25)            <= s_out2(54,26);
	s_locks_lower_in(53,25) <= s_locks_lower_out(54,25);

		normal_cell_53_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,26),
			fetch              => s_fetch(53,26),
			data_in            => s_data_in(53,26),
			data_out           => s_data_out(53,26),
			out1               => s_out1(53,26),
			out2               => s_out2(53,26),
			lock_lower_row_out => s_locks_lower_out(53,26),
			lock_lower_row_in  => s_locks_lower_in(53,26),
			in1                => s_in1(53,26),
			in2                => s_in2(53,26),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(26)
		);
	s_in1(53,26)            <= s_out1(54,26);
	s_in2(53,26)            <= s_out2(54,27);
	s_locks_lower_in(53,26) <= s_locks_lower_out(54,26);

		normal_cell_53_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,27),
			fetch              => s_fetch(53,27),
			data_in            => s_data_in(53,27),
			data_out           => s_data_out(53,27),
			out1               => s_out1(53,27),
			out2               => s_out2(53,27),
			lock_lower_row_out => s_locks_lower_out(53,27),
			lock_lower_row_in  => s_locks_lower_in(53,27),
			in1                => s_in1(53,27),
			in2                => s_in2(53,27),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(27)
		);
	s_in1(53,27)            <= s_out1(54,27);
	s_in2(53,27)            <= s_out2(54,28);
	s_locks_lower_in(53,27) <= s_locks_lower_out(54,27);

		normal_cell_53_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,28),
			fetch              => s_fetch(53,28),
			data_in            => s_data_in(53,28),
			data_out           => s_data_out(53,28),
			out1               => s_out1(53,28),
			out2               => s_out2(53,28),
			lock_lower_row_out => s_locks_lower_out(53,28),
			lock_lower_row_in  => s_locks_lower_in(53,28),
			in1                => s_in1(53,28),
			in2                => s_in2(53,28),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(28)
		);
	s_in1(53,28)            <= s_out1(54,28);
	s_in2(53,28)            <= s_out2(54,29);
	s_locks_lower_in(53,28) <= s_locks_lower_out(54,28);

		normal_cell_53_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,29),
			fetch              => s_fetch(53,29),
			data_in            => s_data_in(53,29),
			data_out           => s_data_out(53,29),
			out1               => s_out1(53,29),
			out2               => s_out2(53,29),
			lock_lower_row_out => s_locks_lower_out(53,29),
			lock_lower_row_in  => s_locks_lower_in(53,29),
			in1                => s_in1(53,29),
			in2                => s_in2(53,29),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(29)
		);
	s_in1(53,29)            <= s_out1(54,29);
	s_in2(53,29)            <= s_out2(54,30);
	s_locks_lower_in(53,29) <= s_locks_lower_out(54,29);

		normal_cell_53_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,30),
			fetch              => s_fetch(53,30),
			data_in            => s_data_in(53,30),
			data_out           => s_data_out(53,30),
			out1               => s_out1(53,30),
			out2               => s_out2(53,30),
			lock_lower_row_out => s_locks_lower_out(53,30),
			lock_lower_row_in  => s_locks_lower_in(53,30),
			in1                => s_in1(53,30),
			in2                => s_in2(53,30),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(30)
		);
	s_in1(53,30)            <= s_out1(54,30);
	s_in2(53,30)            <= s_out2(54,31);
	s_locks_lower_in(53,30) <= s_locks_lower_out(54,30);

		normal_cell_53_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,31),
			fetch              => s_fetch(53,31),
			data_in            => s_data_in(53,31),
			data_out           => s_data_out(53,31),
			out1               => s_out1(53,31),
			out2               => s_out2(53,31),
			lock_lower_row_out => s_locks_lower_out(53,31),
			lock_lower_row_in  => s_locks_lower_in(53,31),
			in1                => s_in1(53,31),
			in2                => s_in2(53,31),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(31)
		);
	s_in1(53,31)            <= s_out1(54,31);
	s_in2(53,31)            <= s_out2(54,32);
	s_locks_lower_in(53,31) <= s_locks_lower_out(54,31);

		normal_cell_53_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,32),
			fetch              => s_fetch(53,32),
			data_in            => s_data_in(53,32),
			data_out           => s_data_out(53,32),
			out1               => s_out1(53,32),
			out2               => s_out2(53,32),
			lock_lower_row_out => s_locks_lower_out(53,32),
			lock_lower_row_in  => s_locks_lower_in(53,32),
			in1                => s_in1(53,32),
			in2                => s_in2(53,32),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(32)
		);
	s_in1(53,32)            <= s_out1(54,32);
	s_in2(53,32)            <= s_out2(54,33);
	s_locks_lower_in(53,32) <= s_locks_lower_out(54,32);

		normal_cell_53_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,33),
			fetch              => s_fetch(53,33),
			data_in            => s_data_in(53,33),
			data_out           => s_data_out(53,33),
			out1               => s_out1(53,33),
			out2               => s_out2(53,33),
			lock_lower_row_out => s_locks_lower_out(53,33),
			lock_lower_row_in  => s_locks_lower_in(53,33),
			in1                => s_in1(53,33),
			in2                => s_in2(53,33),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(33)
		);
	s_in1(53,33)            <= s_out1(54,33);
	s_in2(53,33)            <= s_out2(54,34);
	s_locks_lower_in(53,33) <= s_locks_lower_out(54,33);

		normal_cell_53_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,34),
			fetch              => s_fetch(53,34),
			data_in            => s_data_in(53,34),
			data_out           => s_data_out(53,34),
			out1               => s_out1(53,34),
			out2               => s_out2(53,34),
			lock_lower_row_out => s_locks_lower_out(53,34),
			lock_lower_row_in  => s_locks_lower_in(53,34),
			in1                => s_in1(53,34),
			in2                => s_in2(53,34),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(34)
		);
	s_in1(53,34)            <= s_out1(54,34);
	s_in2(53,34)            <= s_out2(54,35);
	s_locks_lower_in(53,34) <= s_locks_lower_out(54,34);

		normal_cell_53_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,35),
			fetch              => s_fetch(53,35),
			data_in            => s_data_in(53,35),
			data_out           => s_data_out(53,35),
			out1               => s_out1(53,35),
			out2               => s_out2(53,35),
			lock_lower_row_out => s_locks_lower_out(53,35),
			lock_lower_row_in  => s_locks_lower_in(53,35),
			in1                => s_in1(53,35),
			in2                => s_in2(53,35),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(35)
		);
	s_in1(53,35)            <= s_out1(54,35);
	s_in2(53,35)            <= s_out2(54,36);
	s_locks_lower_in(53,35) <= s_locks_lower_out(54,35);

		normal_cell_53_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,36),
			fetch              => s_fetch(53,36),
			data_in            => s_data_in(53,36),
			data_out           => s_data_out(53,36),
			out1               => s_out1(53,36),
			out2               => s_out2(53,36),
			lock_lower_row_out => s_locks_lower_out(53,36),
			lock_lower_row_in  => s_locks_lower_in(53,36),
			in1                => s_in1(53,36),
			in2                => s_in2(53,36),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(36)
		);
	s_in1(53,36)            <= s_out1(54,36);
	s_in2(53,36)            <= s_out2(54,37);
	s_locks_lower_in(53,36) <= s_locks_lower_out(54,36);

		normal_cell_53_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,37),
			fetch              => s_fetch(53,37),
			data_in            => s_data_in(53,37),
			data_out           => s_data_out(53,37),
			out1               => s_out1(53,37),
			out2               => s_out2(53,37),
			lock_lower_row_out => s_locks_lower_out(53,37),
			lock_lower_row_in  => s_locks_lower_in(53,37),
			in1                => s_in1(53,37),
			in2                => s_in2(53,37),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(37)
		);
	s_in1(53,37)            <= s_out1(54,37);
	s_in2(53,37)            <= s_out2(54,38);
	s_locks_lower_in(53,37) <= s_locks_lower_out(54,37);

		normal_cell_53_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,38),
			fetch              => s_fetch(53,38),
			data_in            => s_data_in(53,38),
			data_out           => s_data_out(53,38),
			out1               => s_out1(53,38),
			out2               => s_out2(53,38),
			lock_lower_row_out => s_locks_lower_out(53,38),
			lock_lower_row_in  => s_locks_lower_in(53,38),
			in1                => s_in1(53,38),
			in2                => s_in2(53,38),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(38)
		);
	s_in1(53,38)            <= s_out1(54,38);
	s_in2(53,38)            <= s_out2(54,39);
	s_locks_lower_in(53,38) <= s_locks_lower_out(54,38);

		normal_cell_53_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,39),
			fetch              => s_fetch(53,39),
			data_in            => s_data_in(53,39),
			data_out           => s_data_out(53,39),
			out1               => s_out1(53,39),
			out2               => s_out2(53,39),
			lock_lower_row_out => s_locks_lower_out(53,39),
			lock_lower_row_in  => s_locks_lower_in(53,39),
			in1                => s_in1(53,39),
			in2                => s_in2(53,39),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(39)
		);
	s_in1(53,39)            <= s_out1(54,39);
	s_in2(53,39)            <= s_out2(54,40);
	s_locks_lower_in(53,39) <= s_locks_lower_out(54,39);

		normal_cell_53_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,40),
			fetch              => s_fetch(53,40),
			data_in            => s_data_in(53,40),
			data_out           => s_data_out(53,40),
			out1               => s_out1(53,40),
			out2               => s_out2(53,40),
			lock_lower_row_out => s_locks_lower_out(53,40),
			lock_lower_row_in  => s_locks_lower_in(53,40),
			in1                => s_in1(53,40),
			in2                => s_in2(53,40),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(40)
		);
	s_in1(53,40)            <= s_out1(54,40);
	s_in2(53,40)            <= s_out2(54,41);
	s_locks_lower_in(53,40) <= s_locks_lower_out(54,40);

		normal_cell_53_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,41),
			fetch              => s_fetch(53,41),
			data_in            => s_data_in(53,41),
			data_out           => s_data_out(53,41),
			out1               => s_out1(53,41),
			out2               => s_out2(53,41),
			lock_lower_row_out => s_locks_lower_out(53,41),
			lock_lower_row_in  => s_locks_lower_in(53,41),
			in1                => s_in1(53,41),
			in2                => s_in2(53,41),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(41)
		);
	s_in1(53,41)            <= s_out1(54,41);
	s_in2(53,41)            <= s_out2(54,42);
	s_locks_lower_in(53,41) <= s_locks_lower_out(54,41);

		normal_cell_53_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,42),
			fetch              => s_fetch(53,42),
			data_in            => s_data_in(53,42),
			data_out           => s_data_out(53,42),
			out1               => s_out1(53,42),
			out2               => s_out2(53,42),
			lock_lower_row_out => s_locks_lower_out(53,42),
			lock_lower_row_in  => s_locks_lower_in(53,42),
			in1                => s_in1(53,42),
			in2                => s_in2(53,42),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(42)
		);
	s_in1(53,42)            <= s_out1(54,42);
	s_in2(53,42)            <= s_out2(54,43);
	s_locks_lower_in(53,42) <= s_locks_lower_out(54,42);

		normal_cell_53_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,43),
			fetch              => s_fetch(53,43),
			data_in            => s_data_in(53,43),
			data_out           => s_data_out(53,43),
			out1               => s_out1(53,43),
			out2               => s_out2(53,43),
			lock_lower_row_out => s_locks_lower_out(53,43),
			lock_lower_row_in  => s_locks_lower_in(53,43),
			in1                => s_in1(53,43),
			in2                => s_in2(53,43),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(43)
		);
	s_in1(53,43)            <= s_out1(54,43);
	s_in2(53,43)            <= s_out2(54,44);
	s_locks_lower_in(53,43) <= s_locks_lower_out(54,43);

		normal_cell_53_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,44),
			fetch              => s_fetch(53,44),
			data_in            => s_data_in(53,44),
			data_out           => s_data_out(53,44),
			out1               => s_out1(53,44),
			out2               => s_out2(53,44),
			lock_lower_row_out => s_locks_lower_out(53,44),
			lock_lower_row_in  => s_locks_lower_in(53,44),
			in1                => s_in1(53,44),
			in2                => s_in2(53,44),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(44)
		);
	s_in1(53,44)            <= s_out1(54,44);
	s_in2(53,44)            <= s_out2(54,45);
	s_locks_lower_in(53,44) <= s_locks_lower_out(54,44);

		normal_cell_53_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,45),
			fetch              => s_fetch(53,45),
			data_in            => s_data_in(53,45),
			data_out           => s_data_out(53,45),
			out1               => s_out1(53,45),
			out2               => s_out2(53,45),
			lock_lower_row_out => s_locks_lower_out(53,45),
			lock_lower_row_in  => s_locks_lower_in(53,45),
			in1                => s_in1(53,45),
			in2                => s_in2(53,45),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(45)
		);
	s_in1(53,45)            <= s_out1(54,45);
	s_in2(53,45)            <= s_out2(54,46);
	s_locks_lower_in(53,45) <= s_locks_lower_out(54,45);

		normal_cell_53_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,46),
			fetch              => s_fetch(53,46),
			data_in            => s_data_in(53,46),
			data_out           => s_data_out(53,46),
			out1               => s_out1(53,46),
			out2               => s_out2(53,46),
			lock_lower_row_out => s_locks_lower_out(53,46),
			lock_lower_row_in  => s_locks_lower_in(53,46),
			in1                => s_in1(53,46),
			in2                => s_in2(53,46),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(46)
		);
	s_in1(53,46)            <= s_out1(54,46);
	s_in2(53,46)            <= s_out2(54,47);
	s_locks_lower_in(53,46) <= s_locks_lower_out(54,46);

		normal_cell_53_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,47),
			fetch              => s_fetch(53,47),
			data_in            => s_data_in(53,47),
			data_out           => s_data_out(53,47),
			out1               => s_out1(53,47),
			out2               => s_out2(53,47),
			lock_lower_row_out => s_locks_lower_out(53,47),
			lock_lower_row_in  => s_locks_lower_in(53,47),
			in1                => s_in1(53,47),
			in2                => s_in2(53,47),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(47)
		);
	s_in1(53,47)            <= s_out1(54,47);
	s_in2(53,47)            <= s_out2(54,48);
	s_locks_lower_in(53,47) <= s_locks_lower_out(54,47);

		normal_cell_53_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,48),
			fetch              => s_fetch(53,48),
			data_in            => s_data_in(53,48),
			data_out           => s_data_out(53,48),
			out1               => s_out1(53,48),
			out2               => s_out2(53,48),
			lock_lower_row_out => s_locks_lower_out(53,48),
			lock_lower_row_in  => s_locks_lower_in(53,48),
			in1                => s_in1(53,48),
			in2                => s_in2(53,48),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(48)
		);
	s_in1(53,48)            <= s_out1(54,48);
	s_in2(53,48)            <= s_out2(54,49);
	s_locks_lower_in(53,48) <= s_locks_lower_out(54,48);

		normal_cell_53_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,49),
			fetch              => s_fetch(53,49),
			data_in            => s_data_in(53,49),
			data_out           => s_data_out(53,49),
			out1               => s_out1(53,49),
			out2               => s_out2(53,49),
			lock_lower_row_out => s_locks_lower_out(53,49),
			lock_lower_row_in  => s_locks_lower_in(53,49),
			in1                => s_in1(53,49),
			in2                => s_in2(53,49),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(49)
		);
	s_in1(53,49)            <= s_out1(54,49);
	s_in2(53,49)            <= s_out2(54,50);
	s_locks_lower_in(53,49) <= s_locks_lower_out(54,49);

		normal_cell_53_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,50),
			fetch              => s_fetch(53,50),
			data_in            => s_data_in(53,50),
			data_out           => s_data_out(53,50),
			out1               => s_out1(53,50),
			out2               => s_out2(53,50),
			lock_lower_row_out => s_locks_lower_out(53,50),
			lock_lower_row_in  => s_locks_lower_in(53,50),
			in1                => s_in1(53,50),
			in2                => s_in2(53,50),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(50)
		);
	s_in1(53,50)            <= s_out1(54,50);
	s_in2(53,50)            <= s_out2(54,51);
	s_locks_lower_in(53,50) <= s_locks_lower_out(54,50);

		normal_cell_53_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,51),
			fetch              => s_fetch(53,51),
			data_in            => s_data_in(53,51),
			data_out           => s_data_out(53,51),
			out1               => s_out1(53,51),
			out2               => s_out2(53,51),
			lock_lower_row_out => s_locks_lower_out(53,51),
			lock_lower_row_in  => s_locks_lower_in(53,51),
			in1                => s_in1(53,51),
			in2                => s_in2(53,51),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(51)
		);
	s_in1(53,51)            <= s_out1(54,51);
	s_in2(53,51)            <= s_out2(54,52);
	s_locks_lower_in(53,51) <= s_locks_lower_out(54,51);

		normal_cell_53_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,52),
			fetch              => s_fetch(53,52),
			data_in            => s_data_in(53,52),
			data_out           => s_data_out(53,52),
			out1               => s_out1(53,52),
			out2               => s_out2(53,52),
			lock_lower_row_out => s_locks_lower_out(53,52),
			lock_lower_row_in  => s_locks_lower_in(53,52),
			in1                => s_in1(53,52),
			in2                => s_in2(53,52),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(52)
		);
	s_in1(53,52)            <= s_out1(54,52);
	s_in2(53,52)            <= s_out2(54,53);
	s_locks_lower_in(53,52) <= s_locks_lower_out(54,52);

		normal_cell_53_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,53),
			fetch              => s_fetch(53,53),
			data_in            => s_data_in(53,53),
			data_out           => s_data_out(53,53),
			out1               => s_out1(53,53),
			out2               => s_out2(53,53),
			lock_lower_row_out => s_locks_lower_out(53,53),
			lock_lower_row_in  => s_locks_lower_in(53,53),
			in1                => s_in1(53,53),
			in2                => s_in2(53,53),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(53)
		);
	s_in1(53,53)            <= s_out1(54,53);
	s_in2(53,53)            <= s_out2(54,54);
	s_locks_lower_in(53,53) <= s_locks_lower_out(54,53);

		normal_cell_53_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,54),
			fetch              => s_fetch(53,54),
			data_in            => s_data_in(53,54),
			data_out           => s_data_out(53,54),
			out1               => s_out1(53,54),
			out2               => s_out2(53,54),
			lock_lower_row_out => s_locks_lower_out(53,54),
			lock_lower_row_in  => s_locks_lower_in(53,54),
			in1                => s_in1(53,54),
			in2                => s_in2(53,54),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(54)
		);
	s_in1(53,54)            <= s_out1(54,54);
	s_in2(53,54)            <= s_out2(54,55);
	s_locks_lower_in(53,54) <= s_locks_lower_out(54,54);

		normal_cell_53_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,55),
			fetch              => s_fetch(53,55),
			data_in            => s_data_in(53,55),
			data_out           => s_data_out(53,55),
			out1               => s_out1(53,55),
			out2               => s_out2(53,55),
			lock_lower_row_out => s_locks_lower_out(53,55),
			lock_lower_row_in  => s_locks_lower_in(53,55),
			in1                => s_in1(53,55),
			in2                => s_in2(53,55),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(55)
		);
	s_in1(53,55)            <= s_out1(54,55);
	s_in2(53,55)            <= s_out2(54,56);
	s_locks_lower_in(53,55) <= s_locks_lower_out(54,55);

		normal_cell_53_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,56),
			fetch              => s_fetch(53,56),
			data_in            => s_data_in(53,56),
			data_out           => s_data_out(53,56),
			out1               => s_out1(53,56),
			out2               => s_out2(53,56),
			lock_lower_row_out => s_locks_lower_out(53,56),
			lock_lower_row_in  => s_locks_lower_in(53,56),
			in1                => s_in1(53,56),
			in2                => s_in2(53,56),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(56)
		);
	s_in1(53,56)            <= s_out1(54,56);
	s_in2(53,56)            <= s_out2(54,57);
	s_locks_lower_in(53,56) <= s_locks_lower_out(54,56);

		normal_cell_53_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,57),
			fetch              => s_fetch(53,57),
			data_in            => s_data_in(53,57),
			data_out           => s_data_out(53,57),
			out1               => s_out1(53,57),
			out2               => s_out2(53,57),
			lock_lower_row_out => s_locks_lower_out(53,57),
			lock_lower_row_in  => s_locks_lower_in(53,57),
			in1                => s_in1(53,57),
			in2                => s_in2(53,57),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(57)
		);
	s_in1(53,57)            <= s_out1(54,57);
	s_in2(53,57)            <= s_out2(54,58);
	s_locks_lower_in(53,57) <= s_locks_lower_out(54,57);

		normal_cell_53_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,58),
			fetch              => s_fetch(53,58),
			data_in            => s_data_in(53,58),
			data_out           => s_data_out(53,58),
			out1               => s_out1(53,58),
			out2               => s_out2(53,58),
			lock_lower_row_out => s_locks_lower_out(53,58),
			lock_lower_row_in  => s_locks_lower_in(53,58),
			in1                => s_in1(53,58),
			in2                => s_in2(53,58),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(58)
		);
	s_in1(53,58)            <= s_out1(54,58);
	s_in2(53,58)            <= s_out2(54,59);
	s_locks_lower_in(53,58) <= s_locks_lower_out(54,58);

		normal_cell_53_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,59),
			fetch              => s_fetch(53,59),
			data_in            => s_data_in(53,59),
			data_out           => s_data_out(53,59),
			out1               => s_out1(53,59),
			out2               => s_out2(53,59),
			lock_lower_row_out => s_locks_lower_out(53,59),
			lock_lower_row_in  => s_locks_lower_in(53,59),
			in1                => s_in1(53,59),
			in2                => s_in2(53,59),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(59)
		);
	s_in1(53,59)            <= s_out1(54,59);
	s_in2(53,59)            <= s_out2(54,60);
	s_locks_lower_in(53,59) <= s_locks_lower_out(54,59);

		last_col_cell_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(53,60),
			fetch              => s_fetch(53,60),
			data_in            => s_data_in(53,60),
			data_out           => s_data_out(53,60),
			out1               => s_out1(53,60),
			out2               => s_out2(53,60),
			lock_lower_row_out => s_locks_lower_out(53,60),
			lock_lower_row_in  => s_locks_lower_in(53,60),
			in1                => s_in1(53,60),
			in2                => (others => '0'),
			lock_row           => s_locks(53),
			piv_found          => s_piv_found,
			row_data           => s_row_data(53),
			col_data           => s_col_data(60)
		);
	s_in1(53,60)            <= s_out1(54,60);
	s_locks_lower_in(53,60) <= s_locks_lower_out(54,60);

		normal_cell_54_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,1),
			fetch              => s_fetch(54,1),
			data_in            => s_data_in(54,1),
			data_out           => s_data_out(54,1),
			out1               => s_out1(54,1),
			out2               => s_out2(54,1),
			lock_lower_row_out => s_locks_lower_out(54,1),
			lock_lower_row_in  => s_locks_lower_in(54,1),
			in1                => s_in1(54,1),
			in2                => s_in2(54,1),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(1)
		);
	s_in1(54,1)            <= s_out1(55,1);
	s_in2(54,1)            <= s_out2(55,2);
	s_locks_lower_in(54,1) <= s_locks_lower_out(55,1);

		normal_cell_54_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,2),
			fetch              => s_fetch(54,2),
			data_in            => s_data_in(54,2),
			data_out           => s_data_out(54,2),
			out1               => s_out1(54,2),
			out2               => s_out2(54,2),
			lock_lower_row_out => s_locks_lower_out(54,2),
			lock_lower_row_in  => s_locks_lower_in(54,2),
			in1                => s_in1(54,2),
			in2                => s_in2(54,2),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(2)
		);
	s_in1(54,2)            <= s_out1(55,2);
	s_in2(54,2)            <= s_out2(55,3);
	s_locks_lower_in(54,2) <= s_locks_lower_out(55,2);

		normal_cell_54_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,3),
			fetch              => s_fetch(54,3),
			data_in            => s_data_in(54,3),
			data_out           => s_data_out(54,3),
			out1               => s_out1(54,3),
			out2               => s_out2(54,3),
			lock_lower_row_out => s_locks_lower_out(54,3),
			lock_lower_row_in  => s_locks_lower_in(54,3),
			in1                => s_in1(54,3),
			in2                => s_in2(54,3),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(3)
		);
	s_in1(54,3)            <= s_out1(55,3);
	s_in2(54,3)            <= s_out2(55,4);
	s_locks_lower_in(54,3) <= s_locks_lower_out(55,3);

		normal_cell_54_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,4),
			fetch              => s_fetch(54,4),
			data_in            => s_data_in(54,4),
			data_out           => s_data_out(54,4),
			out1               => s_out1(54,4),
			out2               => s_out2(54,4),
			lock_lower_row_out => s_locks_lower_out(54,4),
			lock_lower_row_in  => s_locks_lower_in(54,4),
			in1                => s_in1(54,4),
			in2                => s_in2(54,4),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(4)
		);
	s_in1(54,4)            <= s_out1(55,4);
	s_in2(54,4)            <= s_out2(55,5);
	s_locks_lower_in(54,4) <= s_locks_lower_out(55,4);

		normal_cell_54_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,5),
			fetch              => s_fetch(54,5),
			data_in            => s_data_in(54,5),
			data_out           => s_data_out(54,5),
			out1               => s_out1(54,5),
			out2               => s_out2(54,5),
			lock_lower_row_out => s_locks_lower_out(54,5),
			lock_lower_row_in  => s_locks_lower_in(54,5),
			in1                => s_in1(54,5),
			in2                => s_in2(54,5),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(5)
		);
	s_in1(54,5)            <= s_out1(55,5);
	s_in2(54,5)            <= s_out2(55,6);
	s_locks_lower_in(54,5) <= s_locks_lower_out(55,5);

		normal_cell_54_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,6),
			fetch              => s_fetch(54,6),
			data_in            => s_data_in(54,6),
			data_out           => s_data_out(54,6),
			out1               => s_out1(54,6),
			out2               => s_out2(54,6),
			lock_lower_row_out => s_locks_lower_out(54,6),
			lock_lower_row_in  => s_locks_lower_in(54,6),
			in1                => s_in1(54,6),
			in2                => s_in2(54,6),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(6)
		);
	s_in1(54,6)            <= s_out1(55,6);
	s_in2(54,6)            <= s_out2(55,7);
	s_locks_lower_in(54,6) <= s_locks_lower_out(55,6);

		normal_cell_54_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,7),
			fetch              => s_fetch(54,7),
			data_in            => s_data_in(54,7),
			data_out           => s_data_out(54,7),
			out1               => s_out1(54,7),
			out2               => s_out2(54,7),
			lock_lower_row_out => s_locks_lower_out(54,7),
			lock_lower_row_in  => s_locks_lower_in(54,7),
			in1                => s_in1(54,7),
			in2                => s_in2(54,7),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(7)
		);
	s_in1(54,7)            <= s_out1(55,7);
	s_in2(54,7)            <= s_out2(55,8);
	s_locks_lower_in(54,7) <= s_locks_lower_out(55,7);

		normal_cell_54_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,8),
			fetch              => s_fetch(54,8),
			data_in            => s_data_in(54,8),
			data_out           => s_data_out(54,8),
			out1               => s_out1(54,8),
			out2               => s_out2(54,8),
			lock_lower_row_out => s_locks_lower_out(54,8),
			lock_lower_row_in  => s_locks_lower_in(54,8),
			in1                => s_in1(54,8),
			in2                => s_in2(54,8),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(8)
		);
	s_in1(54,8)            <= s_out1(55,8);
	s_in2(54,8)            <= s_out2(55,9);
	s_locks_lower_in(54,8) <= s_locks_lower_out(55,8);

		normal_cell_54_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,9),
			fetch              => s_fetch(54,9),
			data_in            => s_data_in(54,9),
			data_out           => s_data_out(54,9),
			out1               => s_out1(54,9),
			out2               => s_out2(54,9),
			lock_lower_row_out => s_locks_lower_out(54,9),
			lock_lower_row_in  => s_locks_lower_in(54,9),
			in1                => s_in1(54,9),
			in2                => s_in2(54,9),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(9)
		);
	s_in1(54,9)            <= s_out1(55,9);
	s_in2(54,9)            <= s_out2(55,10);
	s_locks_lower_in(54,9) <= s_locks_lower_out(55,9);

		normal_cell_54_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,10),
			fetch              => s_fetch(54,10),
			data_in            => s_data_in(54,10),
			data_out           => s_data_out(54,10),
			out1               => s_out1(54,10),
			out2               => s_out2(54,10),
			lock_lower_row_out => s_locks_lower_out(54,10),
			lock_lower_row_in  => s_locks_lower_in(54,10),
			in1                => s_in1(54,10),
			in2                => s_in2(54,10),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(10)
		);
	s_in1(54,10)            <= s_out1(55,10);
	s_in2(54,10)            <= s_out2(55,11);
	s_locks_lower_in(54,10) <= s_locks_lower_out(55,10);

		normal_cell_54_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,11),
			fetch              => s_fetch(54,11),
			data_in            => s_data_in(54,11),
			data_out           => s_data_out(54,11),
			out1               => s_out1(54,11),
			out2               => s_out2(54,11),
			lock_lower_row_out => s_locks_lower_out(54,11),
			lock_lower_row_in  => s_locks_lower_in(54,11),
			in1                => s_in1(54,11),
			in2                => s_in2(54,11),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(11)
		);
	s_in1(54,11)            <= s_out1(55,11);
	s_in2(54,11)            <= s_out2(55,12);
	s_locks_lower_in(54,11) <= s_locks_lower_out(55,11);

		normal_cell_54_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,12),
			fetch              => s_fetch(54,12),
			data_in            => s_data_in(54,12),
			data_out           => s_data_out(54,12),
			out1               => s_out1(54,12),
			out2               => s_out2(54,12),
			lock_lower_row_out => s_locks_lower_out(54,12),
			lock_lower_row_in  => s_locks_lower_in(54,12),
			in1                => s_in1(54,12),
			in2                => s_in2(54,12),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(12)
		);
	s_in1(54,12)            <= s_out1(55,12);
	s_in2(54,12)            <= s_out2(55,13);
	s_locks_lower_in(54,12) <= s_locks_lower_out(55,12);

		normal_cell_54_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,13),
			fetch              => s_fetch(54,13),
			data_in            => s_data_in(54,13),
			data_out           => s_data_out(54,13),
			out1               => s_out1(54,13),
			out2               => s_out2(54,13),
			lock_lower_row_out => s_locks_lower_out(54,13),
			lock_lower_row_in  => s_locks_lower_in(54,13),
			in1                => s_in1(54,13),
			in2                => s_in2(54,13),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(13)
		);
	s_in1(54,13)            <= s_out1(55,13);
	s_in2(54,13)            <= s_out2(55,14);
	s_locks_lower_in(54,13) <= s_locks_lower_out(55,13);

		normal_cell_54_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,14),
			fetch              => s_fetch(54,14),
			data_in            => s_data_in(54,14),
			data_out           => s_data_out(54,14),
			out1               => s_out1(54,14),
			out2               => s_out2(54,14),
			lock_lower_row_out => s_locks_lower_out(54,14),
			lock_lower_row_in  => s_locks_lower_in(54,14),
			in1                => s_in1(54,14),
			in2                => s_in2(54,14),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(14)
		);
	s_in1(54,14)            <= s_out1(55,14);
	s_in2(54,14)            <= s_out2(55,15);
	s_locks_lower_in(54,14) <= s_locks_lower_out(55,14);

		normal_cell_54_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,15),
			fetch              => s_fetch(54,15),
			data_in            => s_data_in(54,15),
			data_out           => s_data_out(54,15),
			out1               => s_out1(54,15),
			out2               => s_out2(54,15),
			lock_lower_row_out => s_locks_lower_out(54,15),
			lock_lower_row_in  => s_locks_lower_in(54,15),
			in1                => s_in1(54,15),
			in2                => s_in2(54,15),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(15)
		);
	s_in1(54,15)            <= s_out1(55,15);
	s_in2(54,15)            <= s_out2(55,16);
	s_locks_lower_in(54,15) <= s_locks_lower_out(55,15);

		normal_cell_54_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,16),
			fetch              => s_fetch(54,16),
			data_in            => s_data_in(54,16),
			data_out           => s_data_out(54,16),
			out1               => s_out1(54,16),
			out2               => s_out2(54,16),
			lock_lower_row_out => s_locks_lower_out(54,16),
			lock_lower_row_in  => s_locks_lower_in(54,16),
			in1                => s_in1(54,16),
			in2                => s_in2(54,16),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(16)
		);
	s_in1(54,16)            <= s_out1(55,16);
	s_in2(54,16)            <= s_out2(55,17);
	s_locks_lower_in(54,16) <= s_locks_lower_out(55,16);

		normal_cell_54_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,17),
			fetch              => s_fetch(54,17),
			data_in            => s_data_in(54,17),
			data_out           => s_data_out(54,17),
			out1               => s_out1(54,17),
			out2               => s_out2(54,17),
			lock_lower_row_out => s_locks_lower_out(54,17),
			lock_lower_row_in  => s_locks_lower_in(54,17),
			in1                => s_in1(54,17),
			in2                => s_in2(54,17),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(17)
		);
	s_in1(54,17)            <= s_out1(55,17);
	s_in2(54,17)            <= s_out2(55,18);
	s_locks_lower_in(54,17) <= s_locks_lower_out(55,17);

		normal_cell_54_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,18),
			fetch              => s_fetch(54,18),
			data_in            => s_data_in(54,18),
			data_out           => s_data_out(54,18),
			out1               => s_out1(54,18),
			out2               => s_out2(54,18),
			lock_lower_row_out => s_locks_lower_out(54,18),
			lock_lower_row_in  => s_locks_lower_in(54,18),
			in1                => s_in1(54,18),
			in2                => s_in2(54,18),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(18)
		);
	s_in1(54,18)            <= s_out1(55,18);
	s_in2(54,18)            <= s_out2(55,19);
	s_locks_lower_in(54,18) <= s_locks_lower_out(55,18);

		normal_cell_54_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,19),
			fetch              => s_fetch(54,19),
			data_in            => s_data_in(54,19),
			data_out           => s_data_out(54,19),
			out1               => s_out1(54,19),
			out2               => s_out2(54,19),
			lock_lower_row_out => s_locks_lower_out(54,19),
			lock_lower_row_in  => s_locks_lower_in(54,19),
			in1                => s_in1(54,19),
			in2                => s_in2(54,19),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(19)
		);
	s_in1(54,19)            <= s_out1(55,19);
	s_in2(54,19)            <= s_out2(55,20);
	s_locks_lower_in(54,19) <= s_locks_lower_out(55,19);

		normal_cell_54_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,20),
			fetch              => s_fetch(54,20),
			data_in            => s_data_in(54,20),
			data_out           => s_data_out(54,20),
			out1               => s_out1(54,20),
			out2               => s_out2(54,20),
			lock_lower_row_out => s_locks_lower_out(54,20),
			lock_lower_row_in  => s_locks_lower_in(54,20),
			in1                => s_in1(54,20),
			in2                => s_in2(54,20),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(20)
		);
	s_in1(54,20)            <= s_out1(55,20);
	s_in2(54,20)            <= s_out2(55,21);
	s_locks_lower_in(54,20) <= s_locks_lower_out(55,20);

		normal_cell_54_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,21),
			fetch              => s_fetch(54,21),
			data_in            => s_data_in(54,21),
			data_out           => s_data_out(54,21),
			out1               => s_out1(54,21),
			out2               => s_out2(54,21),
			lock_lower_row_out => s_locks_lower_out(54,21),
			lock_lower_row_in  => s_locks_lower_in(54,21),
			in1                => s_in1(54,21),
			in2                => s_in2(54,21),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(21)
		);
	s_in1(54,21)            <= s_out1(55,21);
	s_in2(54,21)            <= s_out2(55,22);
	s_locks_lower_in(54,21) <= s_locks_lower_out(55,21);

		normal_cell_54_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,22),
			fetch              => s_fetch(54,22),
			data_in            => s_data_in(54,22),
			data_out           => s_data_out(54,22),
			out1               => s_out1(54,22),
			out2               => s_out2(54,22),
			lock_lower_row_out => s_locks_lower_out(54,22),
			lock_lower_row_in  => s_locks_lower_in(54,22),
			in1                => s_in1(54,22),
			in2                => s_in2(54,22),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(22)
		);
	s_in1(54,22)            <= s_out1(55,22);
	s_in2(54,22)            <= s_out2(55,23);
	s_locks_lower_in(54,22) <= s_locks_lower_out(55,22);

		normal_cell_54_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,23),
			fetch              => s_fetch(54,23),
			data_in            => s_data_in(54,23),
			data_out           => s_data_out(54,23),
			out1               => s_out1(54,23),
			out2               => s_out2(54,23),
			lock_lower_row_out => s_locks_lower_out(54,23),
			lock_lower_row_in  => s_locks_lower_in(54,23),
			in1                => s_in1(54,23),
			in2                => s_in2(54,23),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(23)
		);
	s_in1(54,23)            <= s_out1(55,23);
	s_in2(54,23)            <= s_out2(55,24);
	s_locks_lower_in(54,23) <= s_locks_lower_out(55,23);

		normal_cell_54_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,24),
			fetch              => s_fetch(54,24),
			data_in            => s_data_in(54,24),
			data_out           => s_data_out(54,24),
			out1               => s_out1(54,24),
			out2               => s_out2(54,24),
			lock_lower_row_out => s_locks_lower_out(54,24),
			lock_lower_row_in  => s_locks_lower_in(54,24),
			in1                => s_in1(54,24),
			in2                => s_in2(54,24),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(24)
		);
	s_in1(54,24)            <= s_out1(55,24);
	s_in2(54,24)            <= s_out2(55,25);
	s_locks_lower_in(54,24) <= s_locks_lower_out(55,24);

		normal_cell_54_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,25),
			fetch              => s_fetch(54,25),
			data_in            => s_data_in(54,25),
			data_out           => s_data_out(54,25),
			out1               => s_out1(54,25),
			out2               => s_out2(54,25),
			lock_lower_row_out => s_locks_lower_out(54,25),
			lock_lower_row_in  => s_locks_lower_in(54,25),
			in1                => s_in1(54,25),
			in2                => s_in2(54,25),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(25)
		);
	s_in1(54,25)            <= s_out1(55,25);
	s_in2(54,25)            <= s_out2(55,26);
	s_locks_lower_in(54,25) <= s_locks_lower_out(55,25);

		normal_cell_54_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,26),
			fetch              => s_fetch(54,26),
			data_in            => s_data_in(54,26),
			data_out           => s_data_out(54,26),
			out1               => s_out1(54,26),
			out2               => s_out2(54,26),
			lock_lower_row_out => s_locks_lower_out(54,26),
			lock_lower_row_in  => s_locks_lower_in(54,26),
			in1                => s_in1(54,26),
			in2                => s_in2(54,26),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(26)
		);
	s_in1(54,26)            <= s_out1(55,26);
	s_in2(54,26)            <= s_out2(55,27);
	s_locks_lower_in(54,26) <= s_locks_lower_out(55,26);

		normal_cell_54_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,27),
			fetch              => s_fetch(54,27),
			data_in            => s_data_in(54,27),
			data_out           => s_data_out(54,27),
			out1               => s_out1(54,27),
			out2               => s_out2(54,27),
			lock_lower_row_out => s_locks_lower_out(54,27),
			lock_lower_row_in  => s_locks_lower_in(54,27),
			in1                => s_in1(54,27),
			in2                => s_in2(54,27),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(27)
		);
	s_in1(54,27)            <= s_out1(55,27);
	s_in2(54,27)            <= s_out2(55,28);
	s_locks_lower_in(54,27) <= s_locks_lower_out(55,27);

		normal_cell_54_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,28),
			fetch              => s_fetch(54,28),
			data_in            => s_data_in(54,28),
			data_out           => s_data_out(54,28),
			out1               => s_out1(54,28),
			out2               => s_out2(54,28),
			lock_lower_row_out => s_locks_lower_out(54,28),
			lock_lower_row_in  => s_locks_lower_in(54,28),
			in1                => s_in1(54,28),
			in2                => s_in2(54,28),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(28)
		);
	s_in1(54,28)            <= s_out1(55,28);
	s_in2(54,28)            <= s_out2(55,29);
	s_locks_lower_in(54,28) <= s_locks_lower_out(55,28);

		normal_cell_54_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,29),
			fetch              => s_fetch(54,29),
			data_in            => s_data_in(54,29),
			data_out           => s_data_out(54,29),
			out1               => s_out1(54,29),
			out2               => s_out2(54,29),
			lock_lower_row_out => s_locks_lower_out(54,29),
			lock_lower_row_in  => s_locks_lower_in(54,29),
			in1                => s_in1(54,29),
			in2                => s_in2(54,29),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(29)
		);
	s_in1(54,29)            <= s_out1(55,29);
	s_in2(54,29)            <= s_out2(55,30);
	s_locks_lower_in(54,29) <= s_locks_lower_out(55,29);

		normal_cell_54_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,30),
			fetch              => s_fetch(54,30),
			data_in            => s_data_in(54,30),
			data_out           => s_data_out(54,30),
			out1               => s_out1(54,30),
			out2               => s_out2(54,30),
			lock_lower_row_out => s_locks_lower_out(54,30),
			lock_lower_row_in  => s_locks_lower_in(54,30),
			in1                => s_in1(54,30),
			in2                => s_in2(54,30),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(30)
		);
	s_in1(54,30)            <= s_out1(55,30);
	s_in2(54,30)            <= s_out2(55,31);
	s_locks_lower_in(54,30) <= s_locks_lower_out(55,30);

		normal_cell_54_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,31),
			fetch              => s_fetch(54,31),
			data_in            => s_data_in(54,31),
			data_out           => s_data_out(54,31),
			out1               => s_out1(54,31),
			out2               => s_out2(54,31),
			lock_lower_row_out => s_locks_lower_out(54,31),
			lock_lower_row_in  => s_locks_lower_in(54,31),
			in1                => s_in1(54,31),
			in2                => s_in2(54,31),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(31)
		);
	s_in1(54,31)            <= s_out1(55,31);
	s_in2(54,31)            <= s_out2(55,32);
	s_locks_lower_in(54,31) <= s_locks_lower_out(55,31);

		normal_cell_54_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,32),
			fetch              => s_fetch(54,32),
			data_in            => s_data_in(54,32),
			data_out           => s_data_out(54,32),
			out1               => s_out1(54,32),
			out2               => s_out2(54,32),
			lock_lower_row_out => s_locks_lower_out(54,32),
			lock_lower_row_in  => s_locks_lower_in(54,32),
			in1                => s_in1(54,32),
			in2                => s_in2(54,32),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(32)
		);
	s_in1(54,32)            <= s_out1(55,32);
	s_in2(54,32)            <= s_out2(55,33);
	s_locks_lower_in(54,32) <= s_locks_lower_out(55,32);

		normal_cell_54_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,33),
			fetch              => s_fetch(54,33),
			data_in            => s_data_in(54,33),
			data_out           => s_data_out(54,33),
			out1               => s_out1(54,33),
			out2               => s_out2(54,33),
			lock_lower_row_out => s_locks_lower_out(54,33),
			lock_lower_row_in  => s_locks_lower_in(54,33),
			in1                => s_in1(54,33),
			in2                => s_in2(54,33),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(33)
		);
	s_in1(54,33)            <= s_out1(55,33);
	s_in2(54,33)            <= s_out2(55,34);
	s_locks_lower_in(54,33) <= s_locks_lower_out(55,33);

		normal_cell_54_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,34),
			fetch              => s_fetch(54,34),
			data_in            => s_data_in(54,34),
			data_out           => s_data_out(54,34),
			out1               => s_out1(54,34),
			out2               => s_out2(54,34),
			lock_lower_row_out => s_locks_lower_out(54,34),
			lock_lower_row_in  => s_locks_lower_in(54,34),
			in1                => s_in1(54,34),
			in2                => s_in2(54,34),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(34)
		);
	s_in1(54,34)            <= s_out1(55,34);
	s_in2(54,34)            <= s_out2(55,35);
	s_locks_lower_in(54,34) <= s_locks_lower_out(55,34);

		normal_cell_54_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,35),
			fetch              => s_fetch(54,35),
			data_in            => s_data_in(54,35),
			data_out           => s_data_out(54,35),
			out1               => s_out1(54,35),
			out2               => s_out2(54,35),
			lock_lower_row_out => s_locks_lower_out(54,35),
			lock_lower_row_in  => s_locks_lower_in(54,35),
			in1                => s_in1(54,35),
			in2                => s_in2(54,35),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(35)
		);
	s_in1(54,35)            <= s_out1(55,35);
	s_in2(54,35)            <= s_out2(55,36);
	s_locks_lower_in(54,35) <= s_locks_lower_out(55,35);

		normal_cell_54_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,36),
			fetch              => s_fetch(54,36),
			data_in            => s_data_in(54,36),
			data_out           => s_data_out(54,36),
			out1               => s_out1(54,36),
			out2               => s_out2(54,36),
			lock_lower_row_out => s_locks_lower_out(54,36),
			lock_lower_row_in  => s_locks_lower_in(54,36),
			in1                => s_in1(54,36),
			in2                => s_in2(54,36),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(36)
		);
	s_in1(54,36)            <= s_out1(55,36);
	s_in2(54,36)            <= s_out2(55,37);
	s_locks_lower_in(54,36) <= s_locks_lower_out(55,36);

		normal_cell_54_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,37),
			fetch              => s_fetch(54,37),
			data_in            => s_data_in(54,37),
			data_out           => s_data_out(54,37),
			out1               => s_out1(54,37),
			out2               => s_out2(54,37),
			lock_lower_row_out => s_locks_lower_out(54,37),
			lock_lower_row_in  => s_locks_lower_in(54,37),
			in1                => s_in1(54,37),
			in2                => s_in2(54,37),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(37)
		);
	s_in1(54,37)            <= s_out1(55,37);
	s_in2(54,37)            <= s_out2(55,38);
	s_locks_lower_in(54,37) <= s_locks_lower_out(55,37);

		normal_cell_54_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,38),
			fetch              => s_fetch(54,38),
			data_in            => s_data_in(54,38),
			data_out           => s_data_out(54,38),
			out1               => s_out1(54,38),
			out2               => s_out2(54,38),
			lock_lower_row_out => s_locks_lower_out(54,38),
			lock_lower_row_in  => s_locks_lower_in(54,38),
			in1                => s_in1(54,38),
			in2                => s_in2(54,38),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(38)
		);
	s_in1(54,38)            <= s_out1(55,38);
	s_in2(54,38)            <= s_out2(55,39);
	s_locks_lower_in(54,38) <= s_locks_lower_out(55,38);

		normal_cell_54_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,39),
			fetch              => s_fetch(54,39),
			data_in            => s_data_in(54,39),
			data_out           => s_data_out(54,39),
			out1               => s_out1(54,39),
			out2               => s_out2(54,39),
			lock_lower_row_out => s_locks_lower_out(54,39),
			lock_lower_row_in  => s_locks_lower_in(54,39),
			in1                => s_in1(54,39),
			in2                => s_in2(54,39),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(39)
		);
	s_in1(54,39)            <= s_out1(55,39);
	s_in2(54,39)            <= s_out2(55,40);
	s_locks_lower_in(54,39) <= s_locks_lower_out(55,39);

		normal_cell_54_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,40),
			fetch              => s_fetch(54,40),
			data_in            => s_data_in(54,40),
			data_out           => s_data_out(54,40),
			out1               => s_out1(54,40),
			out2               => s_out2(54,40),
			lock_lower_row_out => s_locks_lower_out(54,40),
			lock_lower_row_in  => s_locks_lower_in(54,40),
			in1                => s_in1(54,40),
			in2                => s_in2(54,40),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(40)
		);
	s_in1(54,40)            <= s_out1(55,40);
	s_in2(54,40)            <= s_out2(55,41);
	s_locks_lower_in(54,40) <= s_locks_lower_out(55,40);

		normal_cell_54_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,41),
			fetch              => s_fetch(54,41),
			data_in            => s_data_in(54,41),
			data_out           => s_data_out(54,41),
			out1               => s_out1(54,41),
			out2               => s_out2(54,41),
			lock_lower_row_out => s_locks_lower_out(54,41),
			lock_lower_row_in  => s_locks_lower_in(54,41),
			in1                => s_in1(54,41),
			in2                => s_in2(54,41),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(41)
		);
	s_in1(54,41)            <= s_out1(55,41);
	s_in2(54,41)            <= s_out2(55,42);
	s_locks_lower_in(54,41) <= s_locks_lower_out(55,41);

		normal_cell_54_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,42),
			fetch              => s_fetch(54,42),
			data_in            => s_data_in(54,42),
			data_out           => s_data_out(54,42),
			out1               => s_out1(54,42),
			out2               => s_out2(54,42),
			lock_lower_row_out => s_locks_lower_out(54,42),
			lock_lower_row_in  => s_locks_lower_in(54,42),
			in1                => s_in1(54,42),
			in2                => s_in2(54,42),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(42)
		);
	s_in1(54,42)            <= s_out1(55,42);
	s_in2(54,42)            <= s_out2(55,43);
	s_locks_lower_in(54,42) <= s_locks_lower_out(55,42);

		normal_cell_54_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,43),
			fetch              => s_fetch(54,43),
			data_in            => s_data_in(54,43),
			data_out           => s_data_out(54,43),
			out1               => s_out1(54,43),
			out2               => s_out2(54,43),
			lock_lower_row_out => s_locks_lower_out(54,43),
			lock_lower_row_in  => s_locks_lower_in(54,43),
			in1                => s_in1(54,43),
			in2                => s_in2(54,43),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(43)
		);
	s_in1(54,43)            <= s_out1(55,43);
	s_in2(54,43)            <= s_out2(55,44);
	s_locks_lower_in(54,43) <= s_locks_lower_out(55,43);

		normal_cell_54_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,44),
			fetch              => s_fetch(54,44),
			data_in            => s_data_in(54,44),
			data_out           => s_data_out(54,44),
			out1               => s_out1(54,44),
			out2               => s_out2(54,44),
			lock_lower_row_out => s_locks_lower_out(54,44),
			lock_lower_row_in  => s_locks_lower_in(54,44),
			in1                => s_in1(54,44),
			in2                => s_in2(54,44),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(44)
		);
	s_in1(54,44)            <= s_out1(55,44);
	s_in2(54,44)            <= s_out2(55,45);
	s_locks_lower_in(54,44) <= s_locks_lower_out(55,44);

		normal_cell_54_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,45),
			fetch              => s_fetch(54,45),
			data_in            => s_data_in(54,45),
			data_out           => s_data_out(54,45),
			out1               => s_out1(54,45),
			out2               => s_out2(54,45),
			lock_lower_row_out => s_locks_lower_out(54,45),
			lock_lower_row_in  => s_locks_lower_in(54,45),
			in1                => s_in1(54,45),
			in2                => s_in2(54,45),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(45)
		);
	s_in1(54,45)            <= s_out1(55,45);
	s_in2(54,45)            <= s_out2(55,46);
	s_locks_lower_in(54,45) <= s_locks_lower_out(55,45);

		normal_cell_54_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,46),
			fetch              => s_fetch(54,46),
			data_in            => s_data_in(54,46),
			data_out           => s_data_out(54,46),
			out1               => s_out1(54,46),
			out2               => s_out2(54,46),
			lock_lower_row_out => s_locks_lower_out(54,46),
			lock_lower_row_in  => s_locks_lower_in(54,46),
			in1                => s_in1(54,46),
			in2                => s_in2(54,46),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(46)
		);
	s_in1(54,46)            <= s_out1(55,46);
	s_in2(54,46)            <= s_out2(55,47);
	s_locks_lower_in(54,46) <= s_locks_lower_out(55,46);

		normal_cell_54_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,47),
			fetch              => s_fetch(54,47),
			data_in            => s_data_in(54,47),
			data_out           => s_data_out(54,47),
			out1               => s_out1(54,47),
			out2               => s_out2(54,47),
			lock_lower_row_out => s_locks_lower_out(54,47),
			lock_lower_row_in  => s_locks_lower_in(54,47),
			in1                => s_in1(54,47),
			in2                => s_in2(54,47),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(47)
		);
	s_in1(54,47)            <= s_out1(55,47);
	s_in2(54,47)            <= s_out2(55,48);
	s_locks_lower_in(54,47) <= s_locks_lower_out(55,47);

		normal_cell_54_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,48),
			fetch              => s_fetch(54,48),
			data_in            => s_data_in(54,48),
			data_out           => s_data_out(54,48),
			out1               => s_out1(54,48),
			out2               => s_out2(54,48),
			lock_lower_row_out => s_locks_lower_out(54,48),
			lock_lower_row_in  => s_locks_lower_in(54,48),
			in1                => s_in1(54,48),
			in2                => s_in2(54,48),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(48)
		);
	s_in1(54,48)            <= s_out1(55,48);
	s_in2(54,48)            <= s_out2(55,49);
	s_locks_lower_in(54,48) <= s_locks_lower_out(55,48);

		normal_cell_54_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,49),
			fetch              => s_fetch(54,49),
			data_in            => s_data_in(54,49),
			data_out           => s_data_out(54,49),
			out1               => s_out1(54,49),
			out2               => s_out2(54,49),
			lock_lower_row_out => s_locks_lower_out(54,49),
			lock_lower_row_in  => s_locks_lower_in(54,49),
			in1                => s_in1(54,49),
			in2                => s_in2(54,49),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(49)
		);
	s_in1(54,49)            <= s_out1(55,49);
	s_in2(54,49)            <= s_out2(55,50);
	s_locks_lower_in(54,49) <= s_locks_lower_out(55,49);

		normal_cell_54_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,50),
			fetch              => s_fetch(54,50),
			data_in            => s_data_in(54,50),
			data_out           => s_data_out(54,50),
			out1               => s_out1(54,50),
			out2               => s_out2(54,50),
			lock_lower_row_out => s_locks_lower_out(54,50),
			lock_lower_row_in  => s_locks_lower_in(54,50),
			in1                => s_in1(54,50),
			in2                => s_in2(54,50),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(50)
		);
	s_in1(54,50)            <= s_out1(55,50);
	s_in2(54,50)            <= s_out2(55,51);
	s_locks_lower_in(54,50) <= s_locks_lower_out(55,50);

		normal_cell_54_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,51),
			fetch              => s_fetch(54,51),
			data_in            => s_data_in(54,51),
			data_out           => s_data_out(54,51),
			out1               => s_out1(54,51),
			out2               => s_out2(54,51),
			lock_lower_row_out => s_locks_lower_out(54,51),
			lock_lower_row_in  => s_locks_lower_in(54,51),
			in1                => s_in1(54,51),
			in2                => s_in2(54,51),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(51)
		);
	s_in1(54,51)            <= s_out1(55,51);
	s_in2(54,51)            <= s_out2(55,52);
	s_locks_lower_in(54,51) <= s_locks_lower_out(55,51);

		normal_cell_54_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,52),
			fetch              => s_fetch(54,52),
			data_in            => s_data_in(54,52),
			data_out           => s_data_out(54,52),
			out1               => s_out1(54,52),
			out2               => s_out2(54,52),
			lock_lower_row_out => s_locks_lower_out(54,52),
			lock_lower_row_in  => s_locks_lower_in(54,52),
			in1                => s_in1(54,52),
			in2                => s_in2(54,52),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(52)
		);
	s_in1(54,52)            <= s_out1(55,52);
	s_in2(54,52)            <= s_out2(55,53);
	s_locks_lower_in(54,52) <= s_locks_lower_out(55,52);

		normal_cell_54_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,53),
			fetch              => s_fetch(54,53),
			data_in            => s_data_in(54,53),
			data_out           => s_data_out(54,53),
			out1               => s_out1(54,53),
			out2               => s_out2(54,53),
			lock_lower_row_out => s_locks_lower_out(54,53),
			lock_lower_row_in  => s_locks_lower_in(54,53),
			in1                => s_in1(54,53),
			in2                => s_in2(54,53),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(53)
		);
	s_in1(54,53)            <= s_out1(55,53);
	s_in2(54,53)            <= s_out2(55,54);
	s_locks_lower_in(54,53) <= s_locks_lower_out(55,53);

		normal_cell_54_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,54),
			fetch              => s_fetch(54,54),
			data_in            => s_data_in(54,54),
			data_out           => s_data_out(54,54),
			out1               => s_out1(54,54),
			out2               => s_out2(54,54),
			lock_lower_row_out => s_locks_lower_out(54,54),
			lock_lower_row_in  => s_locks_lower_in(54,54),
			in1                => s_in1(54,54),
			in2                => s_in2(54,54),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(54)
		);
	s_in1(54,54)            <= s_out1(55,54);
	s_in2(54,54)            <= s_out2(55,55);
	s_locks_lower_in(54,54) <= s_locks_lower_out(55,54);

		normal_cell_54_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,55),
			fetch              => s_fetch(54,55),
			data_in            => s_data_in(54,55),
			data_out           => s_data_out(54,55),
			out1               => s_out1(54,55),
			out2               => s_out2(54,55),
			lock_lower_row_out => s_locks_lower_out(54,55),
			lock_lower_row_in  => s_locks_lower_in(54,55),
			in1                => s_in1(54,55),
			in2                => s_in2(54,55),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(55)
		);
	s_in1(54,55)            <= s_out1(55,55);
	s_in2(54,55)            <= s_out2(55,56);
	s_locks_lower_in(54,55) <= s_locks_lower_out(55,55);

		normal_cell_54_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,56),
			fetch              => s_fetch(54,56),
			data_in            => s_data_in(54,56),
			data_out           => s_data_out(54,56),
			out1               => s_out1(54,56),
			out2               => s_out2(54,56),
			lock_lower_row_out => s_locks_lower_out(54,56),
			lock_lower_row_in  => s_locks_lower_in(54,56),
			in1                => s_in1(54,56),
			in2                => s_in2(54,56),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(56)
		);
	s_in1(54,56)            <= s_out1(55,56);
	s_in2(54,56)            <= s_out2(55,57);
	s_locks_lower_in(54,56) <= s_locks_lower_out(55,56);

		normal_cell_54_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,57),
			fetch              => s_fetch(54,57),
			data_in            => s_data_in(54,57),
			data_out           => s_data_out(54,57),
			out1               => s_out1(54,57),
			out2               => s_out2(54,57),
			lock_lower_row_out => s_locks_lower_out(54,57),
			lock_lower_row_in  => s_locks_lower_in(54,57),
			in1                => s_in1(54,57),
			in2                => s_in2(54,57),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(57)
		);
	s_in1(54,57)            <= s_out1(55,57);
	s_in2(54,57)            <= s_out2(55,58);
	s_locks_lower_in(54,57) <= s_locks_lower_out(55,57);

		normal_cell_54_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,58),
			fetch              => s_fetch(54,58),
			data_in            => s_data_in(54,58),
			data_out           => s_data_out(54,58),
			out1               => s_out1(54,58),
			out2               => s_out2(54,58),
			lock_lower_row_out => s_locks_lower_out(54,58),
			lock_lower_row_in  => s_locks_lower_in(54,58),
			in1                => s_in1(54,58),
			in2                => s_in2(54,58),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(58)
		);
	s_in1(54,58)            <= s_out1(55,58);
	s_in2(54,58)            <= s_out2(55,59);
	s_locks_lower_in(54,58) <= s_locks_lower_out(55,58);

		normal_cell_54_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,59),
			fetch              => s_fetch(54,59),
			data_in            => s_data_in(54,59),
			data_out           => s_data_out(54,59),
			out1               => s_out1(54,59),
			out2               => s_out2(54,59),
			lock_lower_row_out => s_locks_lower_out(54,59),
			lock_lower_row_in  => s_locks_lower_in(54,59),
			in1                => s_in1(54,59),
			in2                => s_in2(54,59),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(59)
		);
	s_in1(54,59)            <= s_out1(55,59);
	s_in2(54,59)            <= s_out2(55,60);
	s_locks_lower_in(54,59) <= s_locks_lower_out(55,59);

		last_col_cell_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(54,60),
			fetch              => s_fetch(54,60),
			data_in            => s_data_in(54,60),
			data_out           => s_data_out(54,60),
			out1               => s_out1(54,60),
			out2               => s_out2(54,60),
			lock_lower_row_out => s_locks_lower_out(54,60),
			lock_lower_row_in  => s_locks_lower_in(54,60),
			in1                => s_in1(54,60),
			in2                => (others => '0'),
			lock_row           => s_locks(54),
			piv_found          => s_piv_found,
			row_data           => s_row_data(54),
			col_data           => s_col_data(60)
		);
	s_in1(54,60)            <= s_out1(55,60);
	s_locks_lower_in(54,60) <= s_locks_lower_out(55,60);

		normal_cell_55_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,1),
			fetch              => s_fetch(55,1),
			data_in            => s_data_in(55,1),
			data_out           => s_data_out(55,1),
			out1               => s_out1(55,1),
			out2               => s_out2(55,1),
			lock_lower_row_out => s_locks_lower_out(55,1),
			lock_lower_row_in  => s_locks_lower_in(55,1),
			in1                => s_in1(55,1),
			in2                => s_in2(55,1),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(1)
		);
	s_in1(55,1)            <= s_out1(56,1);
	s_in2(55,1)            <= s_out2(56,2);
	s_locks_lower_in(55,1) <= s_locks_lower_out(56,1);

		normal_cell_55_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,2),
			fetch              => s_fetch(55,2),
			data_in            => s_data_in(55,2),
			data_out           => s_data_out(55,2),
			out1               => s_out1(55,2),
			out2               => s_out2(55,2),
			lock_lower_row_out => s_locks_lower_out(55,2),
			lock_lower_row_in  => s_locks_lower_in(55,2),
			in1                => s_in1(55,2),
			in2                => s_in2(55,2),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(2)
		);
	s_in1(55,2)            <= s_out1(56,2);
	s_in2(55,2)            <= s_out2(56,3);
	s_locks_lower_in(55,2) <= s_locks_lower_out(56,2);

		normal_cell_55_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,3),
			fetch              => s_fetch(55,3),
			data_in            => s_data_in(55,3),
			data_out           => s_data_out(55,3),
			out1               => s_out1(55,3),
			out2               => s_out2(55,3),
			lock_lower_row_out => s_locks_lower_out(55,3),
			lock_lower_row_in  => s_locks_lower_in(55,3),
			in1                => s_in1(55,3),
			in2                => s_in2(55,3),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(3)
		);
	s_in1(55,3)            <= s_out1(56,3);
	s_in2(55,3)            <= s_out2(56,4);
	s_locks_lower_in(55,3) <= s_locks_lower_out(56,3);

		normal_cell_55_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,4),
			fetch              => s_fetch(55,4),
			data_in            => s_data_in(55,4),
			data_out           => s_data_out(55,4),
			out1               => s_out1(55,4),
			out2               => s_out2(55,4),
			lock_lower_row_out => s_locks_lower_out(55,4),
			lock_lower_row_in  => s_locks_lower_in(55,4),
			in1                => s_in1(55,4),
			in2                => s_in2(55,4),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(4)
		);
	s_in1(55,4)            <= s_out1(56,4);
	s_in2(55,4)            <= s_out2(56,5);
	s_locks_lower_in(55,4) <= s_locks_lower_out(56,4);

		normal_cell_55_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,5),
			fetch              => s_fetch(55,5),
			data_in            => s_data_in(55,5),
			data_out           => s_data_out(55,5),
			out1               => s_out1(55,5),
			out2               => s_out2(55,5),
			lock_lower_row_out => s_locks_lower_out(55,5),
			lock_lower_row_in  => s_locks_lower_in(55,5),
			in1                => s_in1(55,5),
			in2                => s_in2(55,5),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(5)
		);
	s_in1(55,5)            <= s_out1(56,5);
	s_in2(55,5)            <= s_out2(56,6);
	s_locks_lower_in(55,5) <= s_locks_lower_out(56,5);

		normal_cell_55_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,6),
			fetch              => s_fetch(55,6),
			data_in            => s_data_in(55,6),
			data_out           => s_data_out(55,6),
			out1               => s_out1(55,6),
			out2               => s_out2(55,6),
			lock_lower_row_out => s_locks_lower_out(55,6),
			lock_lower_row_in  => s_locks_lower_in(55,6),
			in1                => s_in1(55,6),
			in2                => s_in2(55,6),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(6)
		);
	s_in1(55,6)            <= s_out1(56,6);
	s_in2(55,6)            <= s_out2(56,7);
	s_locks_lower_in(55,6) <= s_locks_lower_out(56,6);

		normal_cell_55_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,7),
			fetch              => s_fetch(55,7),
			data_in            => s_data_in(55,7),
			data_out           => s_data_out(55,7),
			out1               => s_out1(55,7),
			out2               => s_out2(55,7),
			lock_lower_row_out => s_locks_lower_out(55,7),
			lock_lower_row_in  => s_locks_lower_in(55,7),
			in1                => s_in1(55,7),
			in2                => s_in2(55,7),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(7)
		);
	s_in1(55,7)            <= s_out1(56,7);
	s_in2(55,7)            <= s_out2(56,8);
	s_locks_lower_in(55,7) <= s_locks_lower_out(56,7);

		normal_cell_55_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,8),
			fetch              => s_fetch(55,8),
			data_in            => s_data_in(55,8),
			data_out           => s_data_out(55,8),
			out1               => s_out1(55,8),
			out2               => s_out2(55,8),
			lock_lower_row_out => s_locks_lower_out(55,8),
			lock_lower_row_in  => s_locks_lower_in(55,8),
			in1                => s_in1(55,8),
			in2                => s_in2(55,8),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(8)
		);
	s_in1(55,8)            <= s_out1(56,8);
	s_in2(55,8)            <= s_out2(56,9);
	s_locks_lower_in(55,8) <= s_locks_lower_out(56,8);

		normal_cell_55_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,9),
			fetch              => s_fetch(55,9),
			data_in            => s_data_in(55,9),
			data_out           => s_data_out(55,9),
			out1               => s_out1(55,9),
			out2               => s_out2(55,9),
			lock_lower_row_out => s_locks_lower_out(55,9),
			lock_lower_row_in  => s_locks_lower_in(55,9),
			in1                => s_in1(55,9),
			in2                => s_in2(55,9),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(9)
		);
	s_in1(55,9)            <= s_out1(56,9);
	s_in2(55,9)            <= s_out2(56,10);
	s_locks_lower_in(55,9) <= s_locks_lower_out(56,9);

		normal_cell_55_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,10),
			fetch              => s_fetch(55,10),
			data_in            => s_data_in(55,10),
			data_out           => s_data_out(55,10),
			out1               => s_out1(55,10),
			out2               => s_out2(55,10),
			lock_lower_row_out => s_locks_lower_out(55,10),
			lock_lower_row_in  => s_locks_lower_in(55,10),
			in1                => s_in1(55,10),
			in2                => s_in2(55,10),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(10)
		);
	s_in1(55,10)            <= s_out1(56,10);
	s_in2(55,10)            <= s_out2(56,11);
	s_locks_lower_in(55,10) <= s_locks_lower_out(56,10);

		normal_cell_55_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,11),
			fetch              => s_fetch(55,11),
			data_in            => s_data_in(55,11),
			data_out           => s_data_out(55,11),
			out1               => s_out1(55,11),
			out2               => s_out2(55,11),
			lock_lower_row_out => s_locks_lower_out(55,11),
			lock_lower_row_in  => s_locks_lower_in(55,11),
			in1                => s_in1(55,11),
			in2                => s_in2(55,11),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(11)
		);
	s_in1(55,11)            <= s_out1(56,11);
	s_in2(55,11)            <= s_out2(56,12);
	s_locks_lower_in(55,11) <= s_locks_lower_out(56,11);

		normal_cell_55_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,12),
			fetch              => s_fetch(55,12),
			data_in            => s_data_in(55,12),
			data_out           => s_data_out(55,12),
			out1               => s_out1(55,12),
			out2               => s_out2(55,12),
			lock_lower_row_out => s_locks_lower_out(55,12),
			lock_lower_row_in  => s_locks_lower_in(55,12),
			in1                => s_in1(55,12),
			in2                => s_in2(55,12),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(12)
		);
	s_in1(55,12)            <= s_out1(56,12);
	s_in2(55,12)            <= s_out2(56,13);
	s_locks_lower_in(55,12) <= s_locks_lower_out(56,12);

		normal_cell_55_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,13),
			fetch              => s_fetch(55,13),
			data_in            => s_data_in(55,13),
			data_out           => s_data_out(55,13),
			out1               => s_out1(55,13),
			out2               => s_out2(55,13),
			lock_lower_row_out => s_locks_lower_out(55,13),
			lock_lower_row_in  => s_locks_lower_in(55,13),
			in1                => s_in1(55,13),
			in2                => s_in2(55,13),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(13)
		);
	s_in1(55,13)            <= s_out1(56,13);
	s_in2(55,13)            <= s_out2(56,14);
	s_locks_lower_in(55,13) <= s_locks_lower_out(56,13);

		normal_cell_55_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,14),
			fetch              => s_fetch(55,14),
			data_in            => s_data_in(55,14),
			data_out           => s_data_out(55,14),
			out1               => s_out1(55,14),
			out2               => s_out2(55,14),
			lock_lower_row_out => s_locks_lower_out(55,14),
			lock_lower_row_in  => s_locks_lower_in(55,14),
			in1                => s_in1(55,14),
			in2                => s_in2(55,14),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(14)
		);
	s_in1(55,14)            <= s_out1(56,14);
	s_in2(55,14)            <= s_out2(56,15);
	s_locks_lower_in(55,14) <= s_locks_lower_out(56,14);

		normal_cell_55_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,15),
			fetch              => s_fetch(55,15),
			data_in            => s_data_in(55,15),
			data_out           => s_data_out(55,15),
			out1               => s_out1(55,15),
			out2               => s_out2(55,15),
			lock_lower_row_out => s_locks_lower_out(55,15),
			lock_lower_row_in  => s_locks_lower_in(55,15),
			in1                => s_in1(55,15),
			in2                => s_in2(55,15),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(15)
		);
	s_in1(55,15)            <= s_out1(56,15);
	s_in2(55,15)            <= s_out2(56,16);
	s_locks_lower_in(55,15) <= s_locks_lower_out(56,15);

		normal_cell_55_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,16),
			fetch              => s_fetch(55,16),
			data_in            => s_data_in(55,16),
			data_out           => s_data_out(55,16),
			out1               => s_out1(55,16),
			out2               => s_out2(55,16),
			lock_lower_row_out => s_locks_lower_out(55,16),
			lock_lower_row_in  => s_locks_lower_in(55,16),
			in1                => s_in1(55,16),
			in2                => s_in2(55,16),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(16)
		);
	s_in1(55,16)            <= s_out1(56,16);
	s_in2(55,16)            <= s_out2(56,17);
	s_locks_lower_in(55,16) <= s_locks_lower_out(56,16);

		normal_cell_55_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,17),
			fetch              => s_fetch(55,17),
			data_in            => s_data_in(55,17),
			data_out           => s_data_out(55,17),
			out1               => s_out1(55,17),
			out2               => s_out2(55,17),
			lock_lower_row_out => s_locks_lower_out(55,17),
			lock_lower_row_in  => s_locks_lower_in(55,17),
			in1                => s_in1(55,17),
			in2                => s_in2(55,17),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(17)
		);
	s_in1(55,17)            <= s_out1(56,17);
	s_in2(55,17)            <= s_out2(56,18);
	s_locks_lower_in(55,17) <= s_locks_lower_out(56,17);

		normal_cell_55_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,18),
			fetch              => s_fetch(55,18),
			data_in            => s_data_in(55,18),
			data_out           => s_data_out(55,18),
			out1               => s_out1(55,18),
			out2               => s_out2(55,18),
			lock_lower_row_out => s_locks_lower_out(55,18),
			lock_lower_row_in  => s_locks_lower_in(55,18),
			in1                => s_in1(55,18),
			in2                => s_in2(55,18),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(18)
		);
	s_in1(55,18)            <= s_out1(56,18);
	s_in2(55,18)            <= s_out2(56,19);
	s_locks_lower_in(55,18) <= s_locks_lower_out(56,18);

		normal_cell_55_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,19),
			fetch              => s_fetch(55,19),
			data_in            => s_data_in(55,19),
			data_out           => s_data_out(55,19),
			out1               => s_out1(55,19),
			out2               => s_out2(55,19),
			lock_lower_row_out => s_locks_lower_out(55,19),
			lock_lower_row_in  => s_locks_lower_in(55,19),
			in1                => s_in1(55,19),
			in2                => s_in2(55,19),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(19)
		);
	s_in1(55,19)            <= s_out1(56,19);
	s_in2(55,19)            <= s_out2(56,20);
	s_locks_lower_in(55,19) <= s_locks_lower_out(56,19);

		normal_cell_55_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,20),
			fetch              => s_fetch(55,20),
			data_in            => s_data_in(55,20),
			data_out           => s_data_out(55,20),
			out1               => s_out1(55,20),
			out2               => s_out2(55,20),
			lock_lower_row_out => s_locks_lower_out(55,20),
			lock_lower_row_in  => s_locks_lower_in(55,20),
			in1                => s_in1(55,20),
			in2                => s_in2(55,20),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(20)
		);
	s_in1(55,20)            <= s_out1(56,20);
	s_in2(55,20)            <= s_out2(56,21);
	s_locks_lower_in(55,20) <= s_locks_lower_out(56,20);

		normal_cell_55_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,21),
			fetch              => s_fetch(55,21),
			data_in            => s_data_in(55,21),
			data_out           => s_data_out(55,21),
			out1               => s_out1(55,21),
			out2               => s_out2(55,21),
			lock_lower_row_out => s_locks_lower_out(55,21),
			lock_lower_row_in  => s_locks_lower_in(55,21),
			in1                => s_in1(55,21),
			in2                => s_in2(55,21),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(21)
		);
	s_in1(55,21)            <= s_out1(56,21);
	s_in2(55,21)            <= s_out2(56,22);
	s_locks_lower_in(55,21) <= s_locks_lower_out(56,21);

		normal_cell_55_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,22),
			fetch              => s_fetch(55,22),
			data_in            => s_data_in(55,22),
			data_out           => s_data_out(55,22),
			out1               => s_out1(55,22),
			out2               => s_out2(55,22),
			lock_lower_row_out => s_locks_lower_out(55,22),
			lock_lower_row_in  => s_locks_lower_in(55,22),
			in1                => s_in1(55,22),
			in2                => s_in2(55,22),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(22)
		);
	s_in1(55,22)            <= s_out1(56,22);
	s_in2(55,22)            <= s_out2(56,23);
	s_locks_lower_in(55,22) <= s_locks_lower_out(56,22);

		normal_cell_55_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,23),
			fetch              => s_fetch(55,23),
			data_in            => s_data_in(55,23),
			data_out           => s_data_out(55,23),
			out1               => s_out1(55,23),
			out2               => s_out2(55,23),
			lock_lower_row_out => s_locks_lower_out(55,23),
			lock_lower_row_in  => s_locks_lower_in(55,23),
			in1                => s_in1(55,23),
			in2                => s_in2(55,23),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(23)
		);
	s_in1(55,23)            <= s_out1(56,23);
	s_in2(55,23)            <= s_out2(56,24);
	s_locks_lower_in(55,23) <= s_locks_lower_out(56,23);

		normal_cell_55_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,24),
			fetch              => s_fetch(55,24),
			data_in            => s_data_in(55,24),
			data_out           => s_data_out(55,24),
			out1               => s_out1(55,24),
			out2               => s_out2(55,24),
			lock_lower_row_out => s_locks_lower_out(55,24),
			lock_lower_row_in  => s_locks_lower_in(55,24),
			in1                => s_in1(55,24),
			in2                => s_in2(55,24),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(24)
		);
	s_in1(55,24)            <= s_out1(56,24);
	s_in2(55,24)            <= s_out2(56,25);
	s_locks_lower_in(55,24) <= s_locks_lower_out(56,24);

		normal_cell_55_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,25),
			fetch              => s_fetch(55,25),
			data_in            => s_data_in(55,25),
			data_out           => s_data_out(55,25),
			out1               => s_out1(55,25),
			out2               => s_out2(55,25),
			lock_lower_row_out => s_locks_lower_out(55,25),
			lock_lower_row_in  => s_locks_lower_in(55,25),
			in1                => s_in1(55,25),
			in2                => s_in2(55,25),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(25)
		);
	s_in1(55,25)            <= s_out1(56,25);
	s_in2(55,25)            <= s_out2(56,26);
	s_locks_lower_in(55,25) <= s_locks_lower_out(56,25);

		normal_cell_55_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,26),
			fetch              => s_fetch(55,26),
			data_in            => s_data_in(55,26),
			data_out           => s_data_out(55,26),
			out1               => s_out1(55,26),
			out2               => s_out2(55,26),
			lock_lower_row_out => s_locks_lower_out(55,26),
			lock_lower_row_in  => s_locks_lower_in(55,26),
			in1                => s_in1(55,26),
			in2                => s_in2(55,26),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(26)
		);
	s_in1(55,26)            <= s_out1(56,26);
	s_in2(55,26)            <= s_out2(56,27);
	s_locks_lower_in(55,26) <= s_locks_lower_out(56,26);

		normal_cell_55_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,27),
			fetch              => s_fetch(55,27),
			data_in            => s_data_in(55,27),
			data_out           => s_data_out(55,27),
			out1               => s_out1(55,27),
			out2               => s_out2(55,27),
			lock_lower_row_out => s_locks_lower_out(55,27),
			lock_lower_row_in  => s_locks_lower_in(55,27),
			in1                => s_in1(55,27),
			in2                => s_in2(55,27),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(27)
		);
	s_in1(55,27)            <= s_out1(56,27);
	s_in2(55,27)            <= s_out2(56,28);
	s_locks_lower_in(55,27) <= s_locks_lower_out(56,27);

		normal_cell_55_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,28),
			fetch              => s_fetch(55,28),
			data_in            => s_data_in(55,28),
			data_out           => s_data_out(55,28),
			out1               => s_out1(55,28),
			out2               => s_out2(55,28),
			lock_lower_row_out => s_locks_lower_out(55,28),
			lock_lower_row_in  => s_locks_lower_in(55,28),
			in1                => s_in1(55,28),
			in2                => s_in2(55,28),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(28)
		);
	s_in1(55,28)            <= s_out1(56,28);
	s_in2(55,28)            <= s_out2(56,29);
	s_locks_lower_in(55,28) <= s_locks_lower_out(56,28);

		normal_cell_55_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,29),
			fetch              => s_fetch(55,29),
			data_in            => s_data_in(55,29),
			data_out           => s_data_out(55,29),
			out1               => s_out1(55,29),
			out2               => s_out2(55,29),
			lock_lower_row_out => s_locks_lower_out(55,29),
			lock_lower_row_in  => s_locks_lower_in(55,29),
			in1                => s_in1(55,29),
			in2                => s_in2(55,29),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(29)
		);
	s_in1(55,29)            <= s_out1(56,29);
	s_in2(55,29)            <= s_out2(56,30);
	s_locks_lower_in(55,29) <= s_locks_lower_out(56,29);

		normal_cell_55_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,30),
			fetch              => s_fetch(55,30),
			data_in            => s_data_in(55,30),
			data_out           => s_data_out(55,30),
			out1               => s_out1(55,30),
			out2               => s_out2(55,30),
			lock_lower_row_out => s_locks_lower_out(55,30),
			lock_lower_row_in  => s_locks_lower_in(55,30),
			in1                => s_in1(55,30),
			in2                => s_in2(55,30),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(30)
		);
	s_in1(55,30)            <= s_out1(56,30);
	s_in2(55,30)            <= s_out2(56,31);
	s_locks_lower_in(55,30) <= s_locks_lower_out(56,30);

		normal_cell_55_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,31),
			fetch              => s_fetch(55,31),
			data_in            => s_data_in(55,31),
			data_out           => s_data_out(55,31),
			out1               => s_out1(55,31),
			out2               => s_out2(55,31),
			lock_lower_row_out => s_locks_lower_out(55,31),
			lock_lower_row_in  => s_locks_lower_in(55,31),
			in1                => s_in1(55,31),
			in2                => s_in2(55,31),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(31)
		);
	s_in1(55,31)            <= s_out1(56,31);
	s_in2(55,31)            <= s_out2(56,32);
	s_locks_lower_in(55,31) <= s_locks_lower_out(56,31);

		normal_cell_55_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,32),
			fetch              => s_fetch(55,32),
			data_in            => s_data_in(55,32),
			data_out           => s_data_out(55,32),
			out1               => s_out1(55,32),
			out2               => s_out2(55,32),
			lock_lower_row_out => s_locks_lower_out(55,32),
			lock_lower_row_in  => s_locks_lower_in(55,32),
			in1                => s_in1(55,32),
			in2                => s_in2(55,32),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(32)
		);
	s_in1(55,32)            <= s_out1(56,32);
	s_in2(55,32)            <= s_out2(56,33);
	s_locks_lower_in(55,32) <= s_locks_lower_out(56,32);

		normal_cell_55_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,33),
			fetch              => s_fetch(55,33),
			data_in            => s_data_in(55,33),
			data_out           => s_data_out(55,33),
			out1               => s_out1(55,33),
			out2               => s_out2(55,33),
			lock_lower_row_out => s_locks_lower_out(55,33),
			lock_lower_row_in  => s_locks_lower_in(55,33),
			in1                => s_in1(55,33),
			in2                => s_in2(55,33),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(33)
		);
	s_in1(55,33)            <= s_out1(56,33);
	s_in2(55,33)            <= s_out2(56,34);
	s_locks_lower_in(55,33) <= s_locks_lower_out(56,33);

		normal_cell_55_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,34),
			fetch              => s_fetch(55,34),
			data_in            => s_data_in(55,34),
			data_out           => s_data_out(55,34),
			out1               => s_out1(55,34),
			out2               => s_out2(55,34),
			lock_lower_row_out => s_locks_lower_out(55,34),
			lock_lower_row_in  => s_locks_lower_in(55,34),
			in1                => s_in1(55,34),
			in2                => s_in2(55,34),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(34)
		);
	s_in1(55,34)            <= s_out1(56,34);
	s_in2(55,34)            <= s_out2(56,35);
	s_locks_lower_in(55,34) <= s_locks_lower_out(56,34);

		normal_cell_55_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,35),
			fetch              => s_fetch(55,35),
			data_in            => s_data_in(55,35),
			data_out           => s_data_out(55,35),
			out1               => s_out1(55,35),
			out2               => s_out2(55,35),
			lock_lower_row_out => s_locks_lower_out(55,35),
			lock_lower_row_in  => s_locks_lower_in(55,35),
			in1                => s_in1(55,35),
			in2                => s_in2(55,35),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(35)
		);
	s_in1(55,35)            <= s_out1(56,35);
	s_in2(55,35)            <= s_out2(56,36);
	s_locks_lower_in(55,35) <= s_locks_lower_out(56,35);

		normal_cell_55_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,36),
			fetch              => s_fetch(55,36),
			data_in            => s_data_in(55,36),
			data_out           => s_data_out(55,36),
			out1               => s_out1(55,36),
			out2               => s_out2(55,36),
			lock_lower_row_out => s_locks_lower_out(55,36),
			lock_lower_row_in  => s_locks_lower_in(55,36),
			in1                => s_in1(55,36),
			in2                => s_in2(55,36),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(36)
		);
	s_in1(55,36)            <= s_out1(56,36);
	s_in2(55,36)            <= s_out2(56,37);
	s_locks_lower_in(55,36) <= s_locks_lower_out(56,36);

		normal_cell_55_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,37),
			fetch              => s_fetch(55,37),
			data_in            => s_data_in(55,37),
			data_out           => s_data_out(55,37),
			out1               => s_out1(55,37),
			out2               => s_out2(55,37),
			lock_lower_row_out => s_locks_lower_out(55,37),
			lock_lower_row_in  => s_locks_lower_in(55,37),
			in1                => s_in1(55,37),
			in2                => s_in2(55,37),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(37)
		);
	s_in1(55,37)            <= s_out1(56,37);
	s_in2(55,37)            <= s_out2(56,38);
	s_locks_lower_in(55,37) <= s_locks_lower_out(56,37);

		normal_cell_55_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,38),
			fetch              => s_fetch(55,38),
			data_in            => s_data_in(55,38),
			data_out           => s_data_out(55,38),
			out1               => s_out1(55,38),
			out2               => s_out2(55,38),
			lock_lower_row_out => s_locks_lower_out(55,38),
			lock_lower_row_in  => s_locks_lower_in(55,38),
			in1                => s_in1(55,38),
			in2                => s_in2(55,38),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(38)
		);
	s_in1(55,38)            <= s_out1(56,38);
	s_in2(55,38)            <= s_out2(56,39);
	s_locks_lower_in(55,38) <= s_locks_lower_out(56,38);

		normal_cell_55_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,39),
			fetch              => s_fetch(55,39),
			data_in            => s_data_in(55,39),
			data_out           => s_data_out(55,39),
			out1               => s_out1(55,39),
			out2               => s_out2(55,39),
			lock_lower_row_out => s_locks_lower_out(55,39),
			lock_lower_row_in  => s_locks_lower_in(55,39),
			in1                => s_in1(55,39),
			in2                => s_in2(55,39),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(39)
		);
	s_in1(55,39)            <= s_out1(56,39);
	s_in2(55,39)            <= s_out2(56,40);
	s_locks_lower_in(55,39) <= s_locks_lower_out(56,39);

		normal_cell_55_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,40),
			fetch              => s_fetch(55,40),
			data_in            => s_data_in(55,40),
			data_out           => s_data_out(55,40),
			out1               => s_out1(55,40),
			out2               => s_out2(55,40),
			lock_lower_row_out => s_locks_lower_out(55,40),
			lock_lower_row_in  => s_locks_lower_in(55,40),
			in1                => s_in1(55,40),
			in2                => s_in2(55,40),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(40)
		);
	s_in1(55,40)            <= s_out1(56,40);
	s_in2(55,40)            <= s_out2(56,41);
	s_locks_lower_in(55,40) <= s_locks_lower_out(56,40);

		normal_cell_55_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,41),
			fetch              => s_fetch(55,41),
			data_in            => s_data_in(55,41),
			data_out           => s_data_out(55,41),
			out1               => s_out1(55,41),
			out2               => s_out2(55,41),
			lock_lower_row_out => s_locks_lower_out(55,41),
			lock_lower_row_in  => s_locks_lower_in(55,41),
			in1                => s_in1(55,41),
			in2                => s_in2(55,41),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(41)
		);
	s_in1(55,41)            <= s_out1(56,41);
	s_in2(55,41)            <= s_out2(56,42);
	s_locks_lower_in(55,41) <= s_locks_lower_out(56,41);

		normal_cell_55_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,42),
			fetch              => s_fetch(55,42),
			data_in            => s_data_in(55,42),
			data_out           => s_data_out(55,42),
			out1               => s_out1(55,42),
			out2               => s_out2(55,42),
			lock_lower_row_out => s_locks_lower_out(55,42),
			lock_lower_row_in  => s_locks_lower_in(55,42),
			in1                => s_in1(55,42),
			in2                => s_in2(55,42),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(42)
		);
	s_in1(55,42)            <= s_out1(56,42);
	s_in2(55,42)            <= s_out2(56,43);
	s_locks_lower_in(55,42) <= s_locks_lower_out(56,42);

		normal_cell_55_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,43),
			fetch              => s_fetch(55,43),
			data_in            => s_data_in(55,43),
			data_out           => s_data_out(55,43),
			out1               => s_out1(55,43),
			out2               => s_out2(55,43),
			lock_lower_row_out => s_locks_lower_out(55,43),
			lock_lower_row_in  => s_locks_lower_in(55,43),
			in1                => s_in1(55,43),
			in2                => s_in2(55,43),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(43)
		);
	s_in1(55,43)            <= s_out1(56,43);
	s_in2(55,43)            <= s_out2(56,44);
	s_locks_lower_in(55,43) <= s_locks_lower_out(56,43);

		normal_cell_55_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,44),
			fetch              => s_fetch(55,44),
			data_in            => s_data_in(55,44),
			data_out           => s_data_out(55,44),
			out1               => s_out1(55,44),
			out2               => s_out2(55,44),
			lock_lower_row_out => s_locks_lower_out(55,44),
			lock_lower_row_in  => s_locks_lower_in(55,44),
			in1                => s_in1(55,44),
			in2                => s_in2(55,44),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(44)
		);
	s_in1(55,44)            <= s_out1(56,44);
	s_in2(55,44)            <= s_out2(56,45);
	s_locks_lower_in(55,44) <= s_locks_lower_out(56,44);

		normal_cell_55_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,45),
			fetch              => s_fetch(55,45),
			data_in            => s_data_in(55,45),
			data_out           => s_data_out(55,45),
			out1               => s_out1(55,45),
			out2               => s_out2(55,45),
			lock_lower_row_out => s_locks_lower_out(55,45),
			lock_lower_row_in  => s_locks_lower_in(55,45),
			in1                => s_in1(55,45),
			in2                => s_in2(55,45),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(45)
		);
	s_in1(55,45)            <= s_out1(56,45);
	s_in2(55,45)            <= s_out2(56,46);
	s_locks_lower_in(55,45) <= s_locks_lower_out(56,45);

		normal_cell_55_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,46),
			fetch              => s_fetch(55,46),
			data_in            => s_data_in(55,46),
			data_out           => s_data_out(55,46),
			out1               => s_out1(55,46),
			out2               => s_out2(55,46),
			lock_lower_row_out => s_locks_lower_out(55,46),
			lock_lower_row_in  => s_locks_lower_in(55,46),
			in1                => s_in1(55,46),
			in2                => s_in2(55,46),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(46)
		);
	s_in1(55,46)            <= s_out1(56,46);
	s_in2(55,46)            <= s_out2(56,47);
	s_locks_lower_in(55,46) <= s_locks_lower_out(56,46);

		normal_cell_55_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,47),
			fetch              => s_fetch(55,47),
			data_in            => s_data_in(55,47),
			data_out           => s_data_out(55,47),
			out1               => s_out1(55,47),
			out2               => s_out2(55,47),
			lock_lower_row_out => s_locks_lower_out(55,47),
			lock_lower_row_in  => s_locks_lower_in(55,47),
			in1                => s_in1(55,47),
			in2                => s_in2(55,47),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(47)
		);
	s_in1(55,47)            <= s_out1(56,47);
	s_in2(55,47)            <= s_out2(56,48);
	s_locks_lower_in(55,47) <= s_locks_lower_out(56,47);

		normal_cell_55_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,48),
			fetch              => s_fetch(55,48),
			data_in            => s_data_in(55,48),
			data_out           => s_data_out(55,48),
			out1               => s_out1(55,48),
			out2               => s_out2(55,48),
			lock_lower_row_out => s_locks_lower_out(55,48),
			lock_lower_row_in  => s_locks_lower_in(55,48),
			in1                => s_in1(55,48),
			in2                => s_in2(55,48),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(48)
		);
	s_in1(55,48)            <= s_out1(56,48);
	s_in2(55,48)            <= s_out2(56,49);
	s_locks_lower_in(55,48) <= s_locks_lower_out(56,48);

		normal_cell_55_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,49),
			fetch              => s_fetch(55,49),
			data_in            => s_data_in(55,49),
			data_out           => s_data_out(55,49),
			out1               => s_out1(55,49),
			out2               => s_out2(55,49),
			lock_lower_row_out => s_locks_lower_out(55,49),
			lock_lower_row_in  => s_locks_lower_in(55,49),
			in1                => s_in1(55,49),
			in2                => s_in2(55,49),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(49)
		);
	s_in1(55,49)            <= s_out1(56,49);
	s_in2(55,49)            <= s_out2(56,50);
	s_locks_lower_in(55,49) <= s_locks_lower_out(56,49);

		normal_cell_55_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,50),
			fetch              => s_fetch(55,50),
			data_in            => s_data_in(55,50),
			data_out           => s_data_out(55,50),
			out1               => s_out1(55,50),
			out2               => s_out2(55,50),
			lock_lower_row_out => s_locks_lower_out(55,50),
			lock_lower_row_in  => s_locks_lower_in(55,50),
			in1                => s_in1(55,50),
			in2                => s_in2(55,50),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(50)
		);
	s_in1(55,50)            <= s_out1(56,50);
	s_in2(55,50)            <= s_out2(56,51);
	s_locks_lower_in(55,50) <= s_locks_lower_out(56,50);

		normal_cell_55_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,51),
			fetch              => s_fetch(55,51),
			data_in            => s_data_in(55,51),
			data_out           => s_data_out(55,51),
			out1               => s_out1(55,51),
			out2               => s_out2(55,51),
			lock_lower_row_out => s_locks_lower_out(55,51),
			lock_lower_row_in  => s_locks_lower_in(55,51),
			in1                => s_in1(55,51),
			in2                => s_in2(55,51),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(51)
		);
	s_in1(55,51)            <= s_out1(56,51);
	s_in2(55,51)            <= s_out2(56,52);
	s_locks_lower_in(55,51) <= s_locks_lower_out(56,51);

		normal_cell_55_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,52),
			fetch              => s_fetch(55,52),
			data_in            => s_data_in(55,52),
			data_out           => s_data_out(55,52),
			out1               => s_out1(55,52),
			out2               => s_out2(55,52),
			lock_lower_row_out => s_locks_lower_out(55,52),
			lock_lower_row_in  => s_locks_lower_in(55,52),
			in1                => s_in1(55,52),
			in2                => s_in2(55,52),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(52)
		);
	s_in1(55,52)            <= s_out1(56,52);
	s_in2(55,52)            <= s_out2(56,53);
	s_locks_lower_in(55,52) <= s_locks_lower_out(56,52);

		normal_cell_55_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,53),
			fetch              => s_fetch(55,53),
			data_in            => s_data_in(55,53),
			data_out           => s_data_out(55,53),
			out1               => s_out1(55,53),
			out2               => s_out2(55,53),
			lock_lower_row_out => s_locks_lower_out(55,53),
			lock_lower_row_in  => s_locks_lower_in(55,53),
			in1                => s_in1(55,53),
			in2                => s_in2(55,53),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(53)
		);
	s_in1(55,53)            <= s_out1(56,53);
	s_in2(55,53)            <= s_out2(56,54);
	s_locks_lower_in(55,53) <= s_locks_lower_out(56,53);

		normal_cell_55_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,54),
			fetch              => s_fetch(55,54),
			data_in            => s_data_in(55,54),
			data_out           => s_data_out(55,54),
			out1               => s_out1(55,54),
			out2               => s_out2(55,54),
			lock_lower_row_out => s_locks_lower_out(55,54),
			lock_lower_row_in  => s_locks_lower_in(55,54),
			in1                => s_in1(55,54),
			in2                => s_in2(55,54),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(54)
		);
	s_in1(55,54)            <= s_out1(56,54);
	s_in2(55,54)            <= s_out2(56,55);
	s_locks_lower_in(55,54) <= s_locks_lower_out(56,54);

		normal_cell_55_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,55),
			fetch              => s_fetch(55,55),
			data_in            => s_data_in(55,55),
			data_out           => s_data_out(55,55),
			out1               => s_out1(55,55),
			out2               => s_out2(55,55),
			lock_lower_row_out => s_locks_lower_out(55,55),
			lock_lower_row_in  => s_locks_lower_in(55,55),
			in1                => s_in1(55,55),
			in2                => s_in2(55,55),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(55)
		);
	s_in1(55,55)            <= s_out1(56,55);
	s_in2(55,55)            <= s_out2(56,56);
	s_locks_lower_in(55,55) <= s_locks_lower_out(56,55);

		normal_cell_55_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,56),
			fetch              => s_fetch(55,56),
			data_in            => s_data_in(55,56),
			data_out           => s_data_out(55,56),
			out1               => s_out1(55,56),
			out2               => s_out2(55,56),
			lock_lower_row_out => s_locks_lower_out(55,56),
			lock_lower_row_in  => s_locks_lower_in(55,56),
			in1                => s_in1(55,56),
			in2                => s_in2(55,56),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(56)
		);
	s_in1(55,56)            <= s_out1(56,56);
	s_in2(55,56)            <= s_out2(56,57);
	s_locks_lower_in(55,56) <= s_locks_lower_out(56,56);

		normal_cell_55_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,57),
			fetch              => s_fetch(55,57),
			data_in            => s_data_in(55,57),
			data_out           => s_data_out(55,57),
			out1               => s_out1(55,57),
			out2               => s_out2(55,57),
			lock_lower_row_out => s_locks_lower_out(55,57),
			lock_lower_row_in  => s_locks_lower_in(55,57),
			in1                => s_in1(55,57),
			in2                => s_in2(55,57),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(57)
		);
	s_in1(55,57)            <= s_out1(56,57);
	s_in2(55,57)            <= s_out2(56,58);
	s_locks_lower_in(55,57) <= s_locks_lower_out(56,57);

		normal_cell_55_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,58),
			fetch              => s_fetch(55,58),
			data_in            => s_data_in(55,58),
			data_out           => s_data_out(55,58),
			out1               => s_out1(55,58),
			out2               => s_out2(55,58),
			lock_lower_row_out => s_locks_lower_out(55,58),
			lock_lower_row_in  => s_locks_lower_in(55,58),
			in1                => s_in1(55,58),
			in2                => s_in2(55,58),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(58)
		);
	s_in1(55,58)            <= s_out1(56,58);
	s_in2(55,58)            <= s_out2(56,59);
	s_locks_lower_in(55,58) <= s_locks_lower_out(56,58);

		normal_cell_55_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,59),
			fetch              => s_fetch(55,59),
			data_in            => s_data_in(55,59),
			data_out           => s_data_out(55,59),
			out1               => s_out1(55,59),
			out2               => s_out2(55,59),
			lock_lower_row_out => s_locks_lower_out(55,59),
			lock_lower_row_in  => s_locks_lower_in(55,59),
			in1                => s_in1(55,59),
			in2                => s_in2(55,59),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(59)
		);
	s_in1(55,59)            <= s_out1(56,59);
	s_in2(55,59)            <= s_out2(56,60);
	s_locks_lower_in(55,59) <= s_locks_lower_out(56,59);

		last_col_cell_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(55,60),
			fetch              => s_fetch(55,60),
			data_in            => s_data_in(55,60),
			data_out           => s_data_out(55,60),
			out1               => s_out1(55,60),
			out2               => s_out2(55,60),
			lock_lower_row_out => s_locks_lower_out(55,60),
			lock_lower_row_in  => s_locks_lower_in(55,60),
			in1                => s_in1(55,60),
			in2                => (others => '0'),
			lock_row           => s_locks(55),
			piv_found          => s_piv_found,
			row_data           => s_row_data(55),
			col_data           => s_col_data(60)
		);
	s_in1(55,60)            <= s_out1(56,60);
	s_locks_lower_in(55,60) <= s_locks_lower_out(56,60);

		normal_cell_56_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,1),
			fetch              => s_fetch(56,1),
			data_in            => s_data_in(56,1),
			data_out           => s_data_out(56,1),
			out1               => s_out1(56,1),
			out2               => s_out2(56,1),
			lock_lower_row_out => s_locks_lower_out(56,1),
			lock_lower_row_in  => s_locks_lower_in(56,1),
			in1                => s_in1(56,1),
			in2                => s_in2(56,1),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(1)
		);
	s_in1(56,1)            <= s_out1(57,1);
	s_in2(56,1)            <= s_out2(57,2);
	s_locks_lower_in(56,1) <= s_locks_lower_out(57,1);

		normal_cell_56_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,2),
			fetch              => s_fetch(56,2),
			data_in            => s_data_in(56,2),
			data_out           => s_data_out(56,2),
			out1               => s_out1(56,2),
			out2               => s_out2(56,2),
			lock_lower_row_out => s_locks_lower_out(56,2),
			lock_lower_row_in  => s_locks_lower_in(56,2),
			in1                => s_in1(56,2),
			in2                => s_in2(56,2),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(2)
		);
	s_in1(56,2)            <= s_out1(57,2);
	s_in2(56,2)            <= s_out2(57,3);
	s_locks_lower_in(56,2) <= s_locks_lower_out(57,2);

		normal_cell_56_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,3),
			fetch              => s_fetch(56,3),
			data_in            => s_data_in(56,3),
			data_out           => s_data_out(56,3),
			out1               => s_out1(56,3),
			out2               => s_out2(56,3),
			lock_lower_row_out => s_locks_lower_out(56,3),
			lock_lower_row_in  => s_locks_lower_in(56,3),
			in1                => s_in1(56,3),
			in2                => s_in2(56,3),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(3)
		);
	s_in1(56,3)            <= s_out1(57,3);
	s_in2(56,3)            <= s_out2(57,4);
	s_locks_lower_in(56,3) <= s_locks_lower_out(57,3);

		normal_cell_56_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,4),
			fetch              => s_fetch(56,4),
			data_in            => s_data_in(56,4),
			data_out           => s_data_out(56,4),
			out1               => s_out1(56,4),
			out2               => s_out2(56,4),
			lock_lower_row_out => s_locks_lower_out(56,4),
			lock_lower_row_in  => s_locks_lower_in(56,4),
			in1                => s_in1(56,4),
			in2                => s_in2(56,4),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(4)
		);
	s_in1(56,4)            <= s_out1(57,4);
	s_in2(56,4)            <= s_out2(57,5);
	s_locks_lower_in(56,4) <= s_locks_lower_out(57,4);

		normal_cell_56_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,5),
			fetch              => s_fetch(56,5),
			data_in            => s_data_in(56,5),
			data_out           => s_data_out(56,5),
			out1               => s_out1(56,5),
			out2               => s_out2(56,5),
			lock_lower_row_out => s_locks_lower_out(56,5),
			lock_lower_row_in  => s_locks_lower_in(56,5),
			in1                => s_in1(56,5),
			in2                => s_in2(56,5),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(5)
		);
	s_in1(56,5)            <= s_out1(57,5);
	s_in2(56,5)            <= s_out2(57,6);
	s_locks_lower_in(56,5) <= s_locks_lower_out(57,5);

		normal_cell_56_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,6),
			fetch              => s_fetch(56,6),
			data_in            => s_data_in(56,6),
			data_out           => s_data_out(56,6),
			out1               => s_out1(56,6),
			out2               => s_out2(56,6),
			lock_lower_row_out => s_locks_lower_out(56,6),
			lock_lower_row_in  => s_locks_lower_in(56,6),
			in1                => s_in1(56,6),
			in2                => s_in2(56,6),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(6)
		);
	s_in1(56,6)            <= s_out1(57,6);
	s_in2(56,6)            <= s_out2(57,7);
	s_locks_lower_in(56,6) <= s_locks_lower_out(57,6);

		normal_cell_56_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,7),
			fetch              => s_fetch(56,7),
			data_in            => s_data_in(56,7),
			data_out           => s_data_out(56,7),
			out1               => s_out1(56,7),
			out2               => s_out2(56,7),
			lock_lower_row_out => s_locks_lower_out(56,7),
			lock_lower_row_in  => s_locks_lower_in(56,7),
			in1                => s_in1(56,7),
			in2                => s_in2(56,7),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(7)
		);
	s_in1(56,7)            <= s_out1(57,7);
	s_in2(56,7)            <= s_out2(57,8);
	s_locks_lower_in(56,7) <= s_locks_lower_out(57,7);

		normal_cell_56_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,8),
			fetch              => s_fetch(56,8),
			data_in            => s_data_in(56,8),
			data_out           => s_data_out(56,8),
			out1               => s_out1(56,8),
			out2               => s_out2(56,8),
			lock_lower_row_out => s_locks_lower_out(56,8),
			lock_lower_row_in  => s_locks_lower_in(56,8),
			in1                => s_in1(56,8),
			in2                => s_in2(56,8),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(8)
		);
	s_in1(56,8)            <= s_out1(57,8);
	s_in2(56,8)            <= s_out2(57,9);
	s_locks_lower_in(56,8) <= s_locks_lower_out(57,8);

		normal_cell_56_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,9),
			fetch              => s_fetch(56,9),
			data_in            => s_data_in(56,9),
			data_out           => s_data_out(56,9),
			out1               => s_out1(56,9),
			out2               => s_out2(56,9),
			lock_lower_row_out => s_locks_lower_out(56,9),
			lock_lower_row_in  => s_locks_lower_in(56,9),
			in1                => s_in1(56,9),
			in2                => s_in2(56,9),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(9)
		);
	s_in1(56,9)            <= s_out1(57,9);
	s_in2(56,9)            <= s_out2(57,10);
	s_locks_lower_in(56,9) <= s_locks_lower_out(57,9);

		normal_cell_56_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,10),
			fetch              => s_fetch(56,10),
			data_in            => s_data_in(56,10),
			data_out           => s_data_out(56,10),
			out1               => s_out1(56,10),
			out2               => s_out2(56,10),
			lock_lower_row_out => s_locks_lower_out(56,10),
			lock_lower_row_in  => s_locks_lower_in(56,10),
			in1                => s_in1(56,10),
			in2                => s_in2(56,10),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(10)
		);
	s_in1(56,10)            <= s_out1(57,10);
	s_in2(56,10)            <= s_out2(57,11);
	s_locks_lower_in(56,10) <= s_locks_lower_out(57,10);

		normal_cell_56_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,11),
			fetch              => s_fetch(56,11),
			data_in            => s_data_in(56,11),
			data_out           => s_data_out(56,11),
			out1               => s_out1(56,11),
			out2               => s_out2(56,11),
			lock_lower_row_out => s_locks_lower_out(56,11),
			lock_lower_row_in  => s_locks_lower_in(56,11),
			in1                => s_in1(56,11),
			in2                => s_in2(56,11),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(11)
		);
	s_in1(56,11)            <= s_out1(57,11);
	s_in2(56,11)            <= s_out2(57,12);
	s_locks_lower_in(56,11) <= s_locks_lower_out(57,11);

		normal_cell_56_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,12),
			fetch              => s_fetch(56,12),
			data_in            => s_data_in(56,12),
			data_out           => s_data_out(56,12),
			out1               => s_out1(56,12),
			out2               => s_out2(56,12),
			lock_lower_row_out => s_locks_lower_out(56,12),
			lock_lower_row_in  => s_locks_lower_in(56,12),
			in1                => s_in1(56,12),
			in2                => s_in2(56,12),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(12)
		);
	s_in1(56,12)            <= s_out1(57,12);
	s_in2(56,12)            <= s_out2(57,13);
	s_locks_lower_in(56,12) <= s_locks_lower_out(57,12);

		normal_cell_56_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,13),
			fetch              => s_fetch(56,13),
			data_in            => s_data_in(56,13),
			data_out           => s_data_out(56,13),
			out1               => s_out1(56,13),
			out2               => s_out2(56,13),
			lock_lower_row_out => s_locks_lower_out(56,13),
			lock_lower_row_in  => s_locks_lower_in(56,13),
			in1                => s_in1(56,13),
			in2                => s_in2(56,13),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(13)
		);
	s_in1(56,13)            <= s_out1(57,13);
	s_in2(56,13)            <= s_out2(57,14);
	s_locks_lower_in(56,13) <= s_locks_lower_out(57,13);

		normal_cell_56_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,14),
			fetch              => s_fetch(56,14),
			data_in            => s_data_in(56,14),
			data_out           => s_data_out(56,14),
			out1               => s_out1(56,14),
			out2               => s_out2(56,14),
			lock_lower_row_out => s_locks_lower_out(56,14),
			lock_lower_row_in  => s_locks_lower_in(56,14),
			in1                => s_in1(56,14),
			in2                => s_in2(56,14),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(14)
		);
	s_in1(56,14)            <= s_out1(57,14);
	s_in2(56,14)            <= s_out2(57,15);
	s_locks_lower_in(56,14) <= s_locks_lower_out(57,14);

		normal_cell_56_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,15),
			fetch              => s_fetch(56,15),
			data_in            => s_data_in(56,15),
			data_out           => s_data_out(56,15),
			out1               => s_out1(56,15),
			out2               => s_out2(56,15),
			lock_lower_row_out => s_locks_lower_out(56,15),
			lock_lower_row_in  => s_locks_lower_in(56,15),
			in1                => s_in1(56,15),
			in2                => s_in2(56,15),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(15)
		);
	s_in1(56,15)            <= s_out1(57,15);
	s_in2(56,15)            <= s_out2(57,16);
	s_locks_lower_in(56,15) <= s_locks_lower_out(57,15);

		normal_cell_56_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,16),
			fetch              => s_fetch(56,16),
			data_in            => s_data_in(56,16),
			data_out           => s_data_out(56,16),
			out1               => s_out1(56,16),
			out2               => s_out2(56,16),
			lock_lower_row_out => s_locks_lower_out(56,16),
			lock_lower_row_in  => s_locks_lower_in(56,16),
			in1                => s_in1(56,16),
			in2                => s_in2(56,16),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(16)
		);
	s_in1(56,16)            <= s_out1(57,16);
	s_in2(56,16)            <= s_out2(57,17);
	s_locks_lower_in(56,16) <= s_locks_lower_out(57,16);

		normal_cell_56_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,17),
			fetch              => s_fetch(56,17),
			data_in            => s_data_in(56,17),
			data_out           => s_data_out(56,17),
			out1               => s_out1(56,17),
			out2               => s_out2(56,17),
			lock_lower_row_out => s_locks_lower_out(56,17),
			lock_lower_row_in  => s_locks_lower_in(56,17),
			in1                => s_in1(56,17),
			in2                => s_in2(56,17),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(17)
		);
	s_in1(56,17)            <= s_out1(57,17);
	s_in2(56,17)            <= s_out2(57,18);
	s_locks_lower_in(56,17) <= s_locks_lower_out(57,17);

		normal_cell_56_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,18),
			fetch              => s_fetch(56,18),
			data_in            => s_data_in(56,18),
			data_out           => s_data_out(56,18),
			out1               => s_out1(56,18),
			out2               => s_out2(56,18),
			lock_lower_row_out => s_locks_lower_out(56,18),
			lock_lower_row_in  => s_locks_lower_in(56,18),
			in1                => s_in1(56,18),
			in2                => s_in2(56,18),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(18)
		);
	s_in1(56,18)            <= s_out1(57,18);
	s_in2(56,18)            <= s_out2(57,19);
	s_locks_lower_in(56,18) <= s_locks_lower_out(57,18);

		normal_cell_56_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,19),
			fetch              => s_fetch(56,19),
			data_in            => s_data_in(56,19),
			data_out           => s_data_out(56,19),
			out1               => s_out1(56,19),
			out2               => s_out2(56,19),
			lock_lower_row_out => s_locks_lower_out(56,19),
			lock_lower_row_in  => s_locks_lower_in(56,19),
			in1                => s_in1(56,19),
			in2                => s_in2(56,19),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(19)
		);
	s_in1(56,19)            <= s_out1(57,19);
	s_in2(56,19)            <= s_out2(57,20);
	s_locks_lower_in(56,19) <= s_locks_lower_out(57,19);

		normal_cell_56_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,20),
			fetch              => s_fetch(56,20),
			data_in            => s_data_in(56,20),
			data_out           => s_data_out(56,20),
			out1               => s_out1(56,20),
			out2               => s_out2(56,20),
			lock_lower_row_out => s_locks_lower_out(56,20),
			lock_lower_row_in  => s_locks_lower_in(56,20),
			in1                => s_in1(56,20),
			in2                => s_in2(56,20),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(20)
		);
	s_in1(56,20)            <= s_out1(57,20);
	s_in2(56,20)            <= s_out2(57,21);
	s_locks_lower_in(56,20) <= s_locks_lower_out(57,20);

		normal_cell_56_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,21),
			fetch              => s_fetch(56,21),
			data_in            => s_data_in(56,21),
			data_out           => s_data_out(56,21),
			out1               => s_out1(56,21),
			out2               => s_out2(56,21),
			lock_lower_row_out => s_locks_lower_out(56,21),
			lock_lower_row_in  => s_locks_lower_in(56,21),
			in1                => s_in1(56,21),
			in2                => s_in2(56,21),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(21)
		);
	s_in1(56,21)            <= s_out1(57,21);
	s_in2(56,21)            <= s_out2(57,22);
	s_locks_lower_in(56,21) <= s_locks_lower_out(57,21);

		normal_cell_56_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,22),
			fetch              => s_fetch(56,22),
			data_in            => s_data_in(56,22),
			data_out           => s_data_out(56,22),
			out1               => s_out1(56,22),
			out2               => s_out2(56,22),
			lock_lower_row_out => s_locks_lower_out(56,22),
			lock_lower_row_in  => s_locks_lower_in(56,22),
			in1                => s_in1(56,22),
			in2                => s_in2(56,22),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(22)
		);
	s_in1(56,22)            <= s_out1(57,22);
	s_in2(56,22)            <= s_out2(57,23);
	s_locks_lower_in(56,22) <= s_locks_lower_out(57,22);

		normal_cell_56_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,23),
			fetch              => s_fetch(56,23),
			data_in            => s_data_in(56,23),
			data_out           => s_data_out(56,23),
			out1               => s_out1(56,23),
			out2               => s_out2(56,23),
			lock_lower_row_out => s_locks_lower_out(56,23),
			lock_lower_row_in  => s_locks_lower_in(56,23),
			in1                => s_in1(56,23),
			in2                => s_in2(56,23),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(23)
		);
	s_in1(56,23)            <= s_out1(57,23);
	s_in2(56,23)            <= s_out2(57,24);
	s_locks_lower_in(56,23) <= s_locks_lower_out(57,23);

		normal_cell_56_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,24),
			fetch              => s_fetch(56,24),
			data_in            => s_data_in(56,24),
			data_out           => s_data_out(56,24),
			out1               => s_out1(56,24),
			out2               => s_out2(56,24),
			lock_lower_row_out => s_locks_lower_out(56,24),
			lock_lower_row_in  => s_locks_lower_in(56,24),
			in1                => s_in1(56,24),
			in2                => s_in2(56,24),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(24)
		);
	s_in1(56,24)            <= s_out1(57,24);
	s_in2(56,24)            <= s_out2(57,25);
	s_locks_lower_in(56,24) <= s_locks_lower_out(57,24);

		normal_cell_56_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,25),
			fetch              => s_fetch(56,25),
			data_in            => s_data_in(56,25),
			data_out           => s_data_out(56,25),
			out1               => s_out1(56,25),
			out2               => s_out2(56,25),
			lock_lower_row_out => s_locks_lower_out(56,25),
			lock_lower_row_in  => s_locks_lower_in(56,25),
			in1                => s_in1(56,25),
			in2                => s_in2(56,25),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(25)
		);
	s_in1(56,25)            <= s_out1(57,25);
	s_in2(56,25)            <= s_out2(57,26);
	s_locks_lower_in(56,25) <= s_locks_lower_out(57,25);

		normal_cell_56_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,26),
			fetch              => s_fetch(56,26),
			data_in            => s_data_in(56,26),
			data_out           => s_data_out(56,26),
			out1               => s_out1(56,26),
			out2               => s_out2(56,26),
			lock_lower_row_out => s_locks_lower_out(56,26),
			lock_lower_row_in  => s_locks_lower_in(56,26),
			in1                => s_in1(56,26),
			in2                => s_in2(56,26),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(26)
		);
	s_in1(56,26)            <= s_out1(57,26);
	s_in2(56,26)            <= s_out2(57,27);
	s_locks_lower_in(56,26) <= s_locks_lower_out(57,26);

		normal_cell_56_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,27),
			fetch              => s_fetch(56,27),
			data_in            => s_data_in(56,27),
			data_out           => s_data_out(56,27),
			out1               => s_out1(56,27),
			out2               => s_out2(56,27),
			lock_lower_row_out => s_locks_lower_out(56,27),
			lock_lower_row_in  => s_locks_lower_in(56,27),
			in1                => s_in1(56,27),
			in2                => s_in2(56,27),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(27)
		);
	s_in1(56,27)            <= s_out1(57,27);
	s_in2(56,27)            <= s_out2(57,28);
	s_locks_lower_in(56,27) <= s_locks_lower_out(57,27);

		normal_cell_56_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,28),
			fetch              => s_fetch(56,28),
			data_in            => s_data_in(56,28),
			data_out           => s_data_out(56,28),
			out1               => s_out1(56,28),
			out2               => s_out2(56,28),
			lock_lower_row_out => s_locks_lower_out(56,28),
			lock_lower_row_in  => s_locks_lower_in(56,28),
			in1                => s_in1(56,28),
			in2                => s_in2(56,28),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(28)
		);
	s_in1(56,28)            <= s_out1(57,28);
	s_in2(56,28)            <= s_out2(57,29);
	s_locks_lower_in(56,28) <= s_locks_lower_out(57,28);

		normal_cell_56_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,29),
			fetch              => s_fetch(56,29),
			data_in            => s_data_in(56,29),
			data_out           => s_data_out(56,29),
			out1               => s_out1(56,29),
			out2               => s_out2(56,29),
			lock_lower_row_out => s_locks_lower_out(56,29),
			lock_lower_row_in  => s_locks_lower_in(56,29),
			in1                => s_in1(56,29),
			in2                => s_in2(56,29),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(29)
		);
	s_in1(56,29)            <= s_out1(57,29);
	s_in2(56,29)            <= s_out2(57,30);
	s_locks_lower_in(56,29) <= s_locks_lower_out(57,29);

		normal_cell_56_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,30),
			fetch              => s_fetch(56,30),
			data_in            => s_data_in(56,30),
			data_out           => s_data_out(56,30),
			out1               => s_out1(56,30),
			out2               => s_out2(56,30),
			lock_lower_row_out => s_locks_lower_out(56,30),
			lock_lower_row_in  => s_locks_lower_in(56,30),
			in1                => s_in1(56,30),
			in2                => s_in2(56,30),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(30)
		);
	s_in1(56,30)            <= s_out1(57,30);
	s_in2(56,30)            <= s_out2(57,31);
	s_locks_lower_in(56,30) <= s_locks_lower_out(57,30);

		normal_cell_56_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,31),
			fetch              => s_fetch(56,31),
			data_in            => s_data_in(56,31),
			data_out           => s_data_out(56,31),
			out1               => s_out1(56,31),
			out2               => s_out2(56,31),
			lock_lower_row_out => s_locks_lower_out(56,31),
			lock_lower_row_in  => s_locks_lower_in(56,31),
			in1                => s_in1(56,31),
			in2                => s_in2(56,31),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(31)
		);
	s_in1(56,31)            <= s_out1(57,31);
	s_in2(56,31)            <= s_out2(57,32);
	s_locks_lower_in(56,31) <= s_locks_lower_out(57,31);

		normal_cell_56_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,32),
			fetch              => s_fetch(56,32),
			data_in            => s_data_in(56,32),
			data_out           => s_data_out(56,32),
			out1               => s_out1(56,32),
			out2               => s_out2(56,32),
			lock_lower_row_out => s_locks_lower_out(56,32),
			lock_lower_row_in  => s_locks_lower_in(56,32),
			in1                => s_in1(56,32),
			in2                => s_in2(56,32),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(32)
		);
	s_in1(56,32)            <= s_out1(57,32);
	s_in2(56,32)            <= s_out2(57,33);
	s_locks_lower_in(56,32) <= s_locks_lower_out(57,32);

		normal_cell_56_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,33),
			fetch              => s_fetch(56,33),
			data_in            => s_data_in(56,33),
			data_out           => s_data_out(56,33),
			out1               => s_out1(56,33),
			out2               => s_out2(56,33),
			lock_lower_row_out => s_locks_lower_out(56,33),
			lock_lower_row_in  => s_locks_lower_in(56,33),
			in1                => s_in1(56,33),
			in2                => s_in2(56,33),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(33)
		);
	s_in1(56,33)            <= s_out1(57,33);
	s_in2(56,33)            <= s_out2(57,34);
	s_locks_lower_in(56,33) <= s_locks_lower_out(57,33);

		normal_cell_56_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,34),
			fetch              => s_fetch(56,34),
			data_in            => s_data_in(56,34),
			data_out           => s_data_out(56,34),
			out1               => s_out1(56,34),
			out2               => s_out2(56,34),
			lock_lower_row_out => s_locks_lower_out(56,34),
			lock_lower_row_in  => s_locks_lower_in(56,34),
			in1                => s_in1(56,34),
			in2                => s_in2(56,34),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(34)
		);
	s_in1(56,34)            <= s_out1(57,34);
	s_in2(56,34)            <= s_out2(57,35);
	s_locks_lower_in(56,34) <= s_locks_lower_out(57,34);

		normal_cell_56_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,35),
			fetch              => s_fetch(56,35),
			data_in            => s_data_in(56,35),
			data_out           => s_data_out(56,35),
			out1               => s_out1(56,35),
			out2               => s_out2(56,35),
			lock_lower_row_out => s_locks_lower_out(56,35),
			lock_lower_row_in  => s_locks_lower_in(56,35),
			in1                => s_in1(56,35),
			in2                => s_in2(56,35),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(35)
		);
	s_in1(56,35)            <= s_out1(57,35);
	s_in2(56,35)            <= s_out2(57,36);
	s_locks_lower_in(56,35) <= s_locks_lower_out(57,35);

		normal_cell_56_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,36),
			fetch              => s_fetch(56,36),
			data_in            => s_data_in(56,36),
			data_out           => s_data_out(56,36),
			out1               => s_out1(56,36),
			out2               => s_out2(56,36),
			lock_lower_row_out => s_locks_lower_out(56,36),
			lock_lower_row_in  => s_locks_lower_in(56,36),
			in1                => s_in1(56,36),
			in2                => s_in2(56,36),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(36)
		);
	s_in1(56,36)            <= s_out1(57,36);
	s_in2(56,36)            <= s_out2(57,37);
	s_locks_lower_in(56,36) <= s_locks_lower_out(57,36);

		normal_cell_56_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,37),
			fetch              => s_fetch(56,37),
			data_in            => s_data_in(56,37),
			data_out           => s_data_out(56,37),
			out1               => s_out1(56,37),
			out2               => s_out2(56,37),
			lock_lower_row_out => s_locks_lower_out(56,37),
			lock_lower_row_in  => s_locks_lower_in(56,37),
			in1                => s_in1(56,37),
			in2                => s_in2(56,37),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(37)
		);
	s_in1(56,37)            <= s_out1(57,37);
	s_in2(56,37)            <= s_out2(57,38);
	s_locks_lower_in(56,37) <= s_locks_lower_out(57,37);

		normal_cell_56_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,38),
			fetch              => s_fetch(56,38),
			data_in            => s_data_in(56,38),
			data_out           => s_data_out(56,38),
			out1               => s_out1(56,38),
			out2               => s_out2(56,38),
			lock_lower_row_out => s_locks_lower_out(56,38),
			lock_lower_row_in  => s_locks_lower_in(56,38),
			in1                => s_in1(56,38),
			in2                => s_in2(56,38),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(38)
		);
	s_in1(56,38)            <= s_out1(57,38);
	s_in2(56,38)            <= s_out2(57,39);
	s_locks_lower_in(56,38) <= s_locks_lower_out(57,38);

		normal_cell_56_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,39),
			fetch              => s_fetch(56,39),
			data_in            => s_data_in(56,39),
			data_out           => s_data_out(56,39),
			out1               => s_out1(56,39),
			out2               => s_out2(56,39),
			lock_lower_row_out => s_locks_lower_out(56,39),
			lock_lower_row_in  => s_locks_lower_in(56,39),
			in1                => s_in1(56,39),
			in2                => s_in2(56,39),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(39)
		);
	s_in1(56,39)            <= s_out1(57,39);
	s_in2(56,39)            <= s_out2(57,40);
	s_locks_lower_in(56,39) <= s_locks_lower_out(57,39);

		normal_cell_56_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,40),
			fetch              => s_fetch(56,40),
			data_in            => s_data_in(56,40),
			data_out           => s_data_out(56,40),
			out1               => s_out1(56,40),
			out2               => s_out2(56,40),
			lock_lower_row_out => s_locks_lower_out(56,40),
			lock_lower_row_in  => s_locks_lower_in(56,40),
			in1                => s_in1(56,40),
			in2                => s_in2(56,40),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(40)
		);
	s_in1(56,40)            <= s_out1(57,40);
	s_in2(56,40)            <= s_out2(57,41);
	s_locks_lower_in(56,40) <= s_locks_lower_out(57,40);

		normal_cell_56_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,41),
			fetch              => s_fetch(56,41),
			data_in            => s_data_in(56,41),
			data_out           => s_data_out(56,41),
			out1               => s_out1(56,41),
			out2               => s_out2(56,41),
			lock_lower_row_out => s_locks_lower_out(56,41),
			lock_lower_row_in  => s_locks_lower_in(56,41),
			in1                => s_in1(56,41),
			in2                => s_in2(56,41),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(41)
		);
	s_in1(56,41)            <= s_out1(57,41);
	s_in2(56,41)            <= s_out2(57,42);
	s_locks_lower_in(56,41) <= s_locks_lower_out(57,41);

		normal_cell_56_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,42),
			fetch              => s_fetch(56,42),
			data_in            => s_data_in(56,42),
			data_out           => s_data_out(56,42),
			out1               => s_out1(56,42),
			out2               => s_out2(56,42),
			lock_lower_row_out => s_locks_lower_out(56,42),
			lock_lower_row_in  => s_locks_lower_in(56,42),
			in1                => s_in1(56,42),
			in2                => s_in2(56,42),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(42)
		);
	s_in1(56,42)            <= s_out1(57,42);
	s_in2(56,42)            <= s_out2(57,43);
	s_locks_lower_in(56,42) <= s_locks_lower_out(57,42);

		normal_cell_56_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,43),
			fetch              => s_fetch(56,43),
			data_in            => s_data_in(56,43),
			data_out           => s_data_out(56,43),
			out1               => s_out1(56,43),
			out2               => s_out2(56,43),
			lock_lower_row_out => s_locks_lower_out(56,43),
			lock_lower_row_in  => s_locks_lower_in(56,43),
			in1                => s_in1(56,43),
			in2                => s_in2(56,43),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(43)
		);
	s_in1(56,43)            <= s_out1(57,43);
	s_in2(56,43)            <= s_out2(57,44);
	s_locks_lower_in(56,43) <= s_locks_lower_out(57,43);

		normal_cell_56_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,44),
			fetch              => s_fetch(56,44),
			data_in            => s_data_in(56,44),
			data_out           => s_data_out(56,44),
			out1               => s_out1(56,44),
			out2               => s_out2(56,44),
			lock_lower_row_out => s_locks_lower_out(56,44),
			lock_lower_row_in  => s_locks_lower_in(56,44),
			in1                => s_in1(56,44),
			in2                => s_in2(56,44),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(44)
		);
	s_in1(56,44)            <= s_out1(57,44);
	s_in2(56,44)            <= s_out2(57,45);
	s_locks_lower_in(56,44) <= s_locks_lower_out(57,44);

		normal_cell_56_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,45),
			fetch              => s_fetch(56,45),
			data_in            => s_data_in(56,45),
			data_out           => s_data_out(56,45),
			out1               => s_out1(56,45),
			out2               => s_out2(56,45),
			lock_lower_row_out => s_locks_lower_out(56,45),
			lock_lower_row_in  => s_locks_lower_in(56,45),
			in1                => s_in1(56,45),
			in2                => s_in2(56,45),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(45)
		);
	s_in1(56,45)            <= s_out1(57,45);
	s_in2(56,45)            <= s_out2(57,46);
	s_locks_lower_in(56,45) <= s_locks_lower_out(57,45);

		normal_cell_56_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,46),
			fetch              => s_fetch(56,46),
			data_in            => s_data_in(56,46),
			data_out           => s_data_out(56,46),
			out1               => s_out1(56,46),
			out2               => s_out2(56,46),
			lock_lower_row_out => s_locks_lower_out(56,46),
			lock_lower_row_in  => s_locks_lower_in(56,46),
			in1                => s_in1(56,46),
			in2                => s_in2(56,46),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(46)
		);
	s_in1(56,46)            <= s_out1(57,46);
	s_in2(56,46)            <= s_out2(57,47);
	s_locks_lower_in(56,46) <= s_locks_lower_out(57,46);

		normal_cell_56_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,47),
			fetch              => s_fetch(56,47),
			data_in            => s_data_in(56,47),
			data_out           => s_data_out(56,47),
			out1               => s_out1(56,47),
			out2               => s_out2(56,47),
			lock_lower_row_out => s_locks_lower_out(56,47),
			lock_lower_row_in  => s_locks_lower_in(56,47),
			in1                => s_in1(56,47),
			in2                => s_in2(56,47),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(47)
		);
	s_in1(56,47)            <= s_out1(57,47);
	s_in2(56,47)            <= s_out2(57,48);
	s_locks_lower_in(56,47) <= s_locks_lower_out(57,47);

		normal_cell_56_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,48),
			fetch              => s_fetch(56,48),
			data_in            => s_data_in(56,48),
			data_out           => s_data_out(56,48),
			out1               => s_out1(56,48),
			out2               => s_out2(56,48),
			lock_lower_row_out => s_locks_lower_out(56,48),
			lock_lower_row_in  => s_locks_lower_in(56,48),
			in1                => s_in1(56,48),
			in2                => s_in2(56,48),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(48)
		);
	s_in1(56,48)            <= s_out1(57,48);
	s_in2(56,48)            <= s_out2(57,49);
	s_locks_lower_in(56,48) <= s_locks_lower_out(57,48);

		normal_cell_56_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,49),
			fetch              => s_fetch(56,49),
			data_in            => s_data_in(56,49),
			data_out           => s_data_out(56,49),
			out1               => s_out1(56,49),
			out2               => s_out2(56,49),
			lock_lower_row_out => s_locks_lower_out(56,49),
			lock_lower_row_in  => s_locks_lower_in(56,49),
			in1                => s_in1(56,49),
			in2                => s_in2(56,49),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(49)
		);
	s_in1(56,49)            <= s_out1(57,49);
	s_in2(56,49)            <= s_out2(57,50);
	s_locks_lower_in(56,49) <= s_locks_lower_out(57,49);

		normal_cell_56_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,50),
			fetch              => s_fetch(56,50),
			data_in            => s_data_in(56,50),
			data_out           => s_data_out(56,50),
			out1               => s_out1(56,50),
			out2               => s_out2(56,50),
			lock_lower_row_out => s_locks_lower_out(56,50),
			lock_lower_row_in  => s_locks_lower_in(56,50),
			in1                => s_in1(56,50),
			in2                => s_in2(56,50),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(50)
		);
	s_in1(56,50)            <= s_out1(57,50);
	s_in2(56,50)            <= s_out2(57,51);
	s_locks_lower_in(56,50) <= s_locks_lower_out(57,50);

		normal_cell_56_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,51),
			fetch              => s_fetch(56,51),
			data_in            => s_data_in(56,51),
			data_out           => s_data_out(56,51),
			out1               => s_out1(56,51),
			out2               => s_out2(56,51),
			lock_lower_row_out => s_locks_lower_out(56,51),
			lock_lower_row_in  => s_locks_lower_in(56,51),
			in1                => s_in1(56,51),
			in2                => s_in2(56,51),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(51)
		);
	s_in1(56,51)            <= s_out1(57,51);
	s_in2(56,51)            <= s_out2(57,52);
	s_locks_lower_in(56,51) <= s_locks_lower_out(57,51);

		normal_cell_56_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,52),
			fetch              => s_fetch(56,52),
			data_in            => s_data_in(56,52),
			data_out           => s_data_out(56,52),
			out1               => s_out1(56,52),
			out2               => s_out2(56,52),
			lock_lower_row_out => s_locks_lower_out(56,52),
			lock_lower_row_in  => s_locks_lower_in(56,52),
			in1                => s_in1(56,52),
			in2                => s_in2(56,52),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(52)
		);
	s_in1(56,52)            <= s_out1(57,52);
	s_in2(56,52)            <= s_out2(57,53);
	s_locks_lower_in(56,52) <= s_locks_lower_out(57,52);

		normal_cell_56_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,53),
			fetch              => s_fetch(56,53),
			data_in            => s_data_in(56,53),
			data_out           => s_data_out(56,53),
			out1               => s_out1(56,53),
			out2               => s_out2(56,53),
			lock_lower_row_out => s_locks_lower_out(56,53),
			lock_lower_row_in  => s_locks_lower_in(56,53),
			in1                => s_in1(56,53),
			in2                => s_in2(56,53),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(53)
		);
	s_in1(56,53)            <= s_out1(57,53);
	s_in2(56,53)            <= s_out2(57,54);
	s_locks_lower_in(56,53) <= s_locks_lower_out(57,53);

		normal_cell_56_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,54),
			fetch              => s_fetch(56,54),
			data_in            => s_data_in(56,54),
			data_out           => s_data_out(56,54),
			out1               => s_out1(56,54),
			out2               => s_out2(56,54),
			lock_lower_row_out => s_locks_lower_out(56,54),
			lock_lower_row_in  => s_locks_lower_in(56,54),
			in1                => s_in1(56,54),
			in2                => s_in2(56,54),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(54)
		);
	s_in1(56,54)            <= s_out1(57,54);
	s_in2(56,54)            <= s_out2(57,55);
	s_locks_lower_in(56,54) <= s_locks_lower_out(57,54);

		normal_cell_56_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,55),
			fetch              => s_fetch(56,55),
			data_in            => s_data_in(56,55),
			data_out           => s_data_out(56,55),
			out1               => s_out1(56,55),
			out2               => s_out2(56,55),
			lock_lower_row_out => s_locks_lower_out(56,55),
			lock_lower_row_in  => s_locks_lower_in(56,55),
			in1                => s_in1(56,55),
			in2                => s_in2(56,55),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(55)
		);
	s_in1(56,55)            <= s_out1(57,55);
	s_in2(56,55)            <= s_out2(57,56);
	s_locks_lower_in(56,55) <= s_locks_lower_out(57,55);

		normal_cell_56_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,56),
			fetch              => s_fetch(56,56),
			data_in            => s_data_in(56,56),
			data_out           => s_data_out(56,56),
			out1               => s_out1(56,56),
			out2               => s_out2(56,56),
			lock_lower_row_out => s_locks_lower_out(56,56),
			lock_lower_row_in  => s_locks_lower_in(56,56),
			in1                => s_in1(56,56),
			in2                => s_in2(56,56),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(56)
		);
	s_in1(56,56)            <= s_out1(57,56);
	s_in2(56,56)            <= s_out2(57,57);
	s_locks_lower_in(56,56) <= s_locks_lower_out(57,56);

		normal_cell_56_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,57),
			fetch              => s_fetch(56,57),
			data_in            => s_data_in(56,57),
			data_out           => s_data_out(56,57),
			out1               => s_out1(56,57),
			out2               => s_out2(56,57),
			lock_lower_row_out => s_locks_lower_out(56,57),
			lock_lower_row_in  => s_locks_lower_in(56,57),
			in1                => s_in1(56,57),
			in2                => s_in2(56,57),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(57)
		);
	s_in1(56,57)            <= s_out1(57,57);
	s_in2(56,57)            <= s_out2(57,58);
	s_locks_lower_in(56,57) <= s_locks_lower_out(57,57);

		normal_cell_56_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,58),
			fetch              => s_fetch(56,58),
			data_in            => s_data_in(56,58),
			data_out           => s_data_out(56,58),
			out1               => s_out1(56,58),
			out2               => s_out2(56,58),
			lock_lower_row_out => s_locks_lower_out(56,58),
			lock_lower_row_in  => s_locks_lower_in(56,58),
			in1                => s_in1(56,58),
			in2                => s_in2(56,58),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(58)
		);
	s_in1(56,58)            <= s_out1(57,58);
	s_in2(56,58)            <= s_out2(57,59);
	s_locks_lower_in(56,58) <= s_locks_lower_out(57,58);

		normal_cell_56_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,59),
			fetch              => s_fetch(56,59),
			data_in            => s_data_in(56,59),
			data_out           => s_data_out(56,59),
			out1               => s_out1(56,59),
			out2               => s_out2(56,59),
			lock_lower_row_out => s_locks_lower_out(56,59),
			lock_lower_row_in  => s_locks_lower_in(56,59),
			in1                => s_in1(56,59),
			in2                => s_in2(56,59),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(59)
		);
	s_in1(56,59)            <= s_out1(57,59);
	s_in2(56,59)            <= s_out2(57,60);
	s_locks_lower_in(56,59) <= s_locks_lower_out(57,59);

		last_col_cell_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(56,60),
			fetch              => s_fetch(56,60),
			data_in            => s_data_in(56,60),
			data_out           => s_data_out(56,60),
			out1               => s_out1(56,60),
			out2               => s_out2(56,60),
			lock_lower_row_out => s_locks_lower_out(56,60),
			lock_lower_row_in  => s_locks_lower_in(56,60),
			in1                => s_in1(56,60),
			in2                => (others => '0'),
			lock_row           => s_locks(56),
			piv_found          => s_piv_found,
			row_data           => s_row_data(56),
			col_data           => s_col_data(60)
		);
	s_in1(56,60)            <= s_out1(57,60);
	s_locks_lower_in(56,60) <= s_locks_lower_out(57,60);

		normal_cell_57_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,1),
			fetch              => s_fetch(57,1),
			data_in            => s_data_in(57,1),
			data_out           => s_data_out(57,1),
			out1               => s_out1(57,1),
			out2               => s_out2(57,1),
			lock_lower_row_out => s_locks_lower_out(57,1),
			lock_lower_row_in  => s_locks_lower_in(57,1),
			in1                => s_in1(57,1),
			in2                => s_in2(57,1),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(1)
		);
	s_in1(57,1)            <= s_out1(58,1);
	s_in2(57,1)            <= s_out2(58,2);
	s_locks_lower_in(57,1) <= s_locks_lower_out(58,1);

		normal_cell_57_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,2),
			fetch              => s_fetch(57,2),
			data_in            => s_data_in(57,2),
			data_out           => s_data_out(57,2),
			out1               => s_out1(57,2),
			out2               => s_out2(57,2),
			lock_lower_row_out => s_locks_lower_out(57,2),
			lock_lower_row_in  => s_locks_lower_in(57,2),
			in1                => s_in1(57,2),
			in2                => s_in2(57,2),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(2)
		);
	s_in1(57,2)            <= s_out1(58,2);
	s_in2(57,2)            <= s_out2(58,3);
	s_locks_lower_in(57,2) <= s_locks_lower_out(58,2);

		normal_cell_57_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,3),
			fetch              => s_fetch(57,3),
			data_in            => s_data_in(57,3),
			data_out           => s_data_out(57,3),
			out1               => s_out1(57,3),
			out2               => s_out2(57,3),
			lock_lower_row_out => s_locks_lower_out(57,3),
			lock_lower_row_in  => s_locks_lower_in(57,3),
			in1                => s_in1(57,3),
			in2                => s_in2(57,3),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(3)
		);
	s_in1(57,3)            <= s_out1(58,3);
	s_in2(57,3)            <= s_out2(58,4);
	s_locks_lower_in(57,3) <= s_locks_lower_out(58,3);

		normal_cell_57_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,4),
			fetch              => s_fetch(57,4),
			data_in            => s_data_in(57,4),
			data_out           => s_data_out(57,4),
			out1               => s_out1(57,4),
			out2               => s_out2(57,4),
			lock_lower_row_out => s_locks_lower_out(57,4),
			lock_lower_row_in  => s_locks_lower_in(57,4),
			in1                => s_in1(57,4),
			in2                => s_in2(57,4),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(4)
		);
	s_in1(57,4)            <= s_out1(58,4);
	s_in2(57,4)            <= s_out2(58,5);
	s_locks_lower_in(57,4) <= s_locks_lower_out(58,4);

		normal_cell_57_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,5),
			fetch              => s_fetch(57,5),
			data_in            => s_data_in(57,5),
			data_out           => s_data_out(57,5),
			out1               => s_out1(57,5),
			out2               => s_out2(57,5),
			lock_lower_row_out => s_locks_lower_out(57,5),
			lock_lower_row_in  => s_locks_lower_in(57,5),
			in1                => s_in1(57,5),
			in2                => s_in2(57,5),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(5)
		);
	s_in1(57,5)            <= s_out1(58,5);
	s_in2(57,5)            <= s_out2(58,6);
	s_locks_lower_in(57,5) <= s_locks_lower_out(58,5);

		normal_cell_57_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,6),
			fetch              => s_fetch(57,6),
			data_in            => s_data_in(57,6),
			data_out           => s_data_out(57,6),
			out1               => s_out1(57,6),
			out2               => s_out2(57,6),
			lock_lower_row_out => s_locks_lower_out(57,6),
			lock_lower_row_in  => s_locks_lower_in(57,6),
			in1                => s_in1(57,6),
			in2                => s_in2(57,6),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(6)
		);
	s_in1(57,6)            <= s_out1(58,6);
	s_in2(57,6)            <= s_out2(58,7);
	s_locks_lower_in(57,6) <= s_locks_lower_out(58,6);

		normal_cell_57_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,7),
			fetch              => s_fetch(57,7),
			data_in            => s_data_in(57,7),
			data_out           => s_data_out(57,7),
			out1               => s_out1(57,7),
			out2               => s_out2(57,7),
			lock_lower_row_out => s_locks_lower_out(57,7),
			lock_lower_row_in  => s_locks_lower_in(57,7),
			in1                => s_in1(57,7),
			in2                => s_in2(57,7),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(7)
		);
	s_in1(57,7)            <= s_out1(58,7);
	s_in2(57,7)            <= s_out2(58,8);
	s_locks_lower_in(57,7) <= s_locks_lower_out(58,7);

		normal_cell_57_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,8),
			fetch              => s_fetch(57,8),
			data_in            => s_data_in(57,8),
			data_out           => s_data_out(57,8),
			out1               => s_out1(57,8),
			out2               => s_out2(57,8),
			lock_lower_row_out => s_locks_lower_out(57,8),
			lock_lower_row_in  => s_locks_lower_in(57,8),
			in1                => s_in1(57,8),
			in2                => s_in2(57,8),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(8)
		);
	s_in1(57,8)            <= s_out1(58,8);
	s_in2(57,8)            <= s_out2(58,9);
	s_locks_lower_in(57,8) <= s_locks_lower_out(58,8);

		normal_cell_57_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,9),
			fetch              => s_fetch(57,9),
			data_in            => s_data_in(57,9),
			data_out           => s_data_out(57,9),
			out1               => s_out1(57,9),
			out2               => s_out2(57,9),
			lock_lower_row_out => s_locks_lower_out(57,9),
			lock_lower_row_in  => s_locks_lower_in(57,9),
			in1                => s_in1(57,9),
			in2                => s_in2(57,9),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(9)
		);
	s_in1(57,9)            <= s_out1(58,9);
	s_in2(57,9)            <= s_out2(58,10);
	s_locks_lower_in(57,9) <= s_locks_lower_out(58,9);

		normal_cell_57_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,10),
			fetch              => s_fetch(57,10),
			data_in            => s_data_in(57,10),
			data_out           => s_data_out(57,10),
			out1               => s_out1(57,10),
			out2               => s_out2(57,10),
			lock_lower_row_out => s_locks_lower_out(57,10),
			lock_lower_row_in  => s_locks_lower_in(57,10),
			in1                => s_in1(57,10),
			in2                => s_in2(57,10),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(10)
		);
	s_in1(57,10)            <= s_out1(58,10);
	s_in2(57,10)            <= s_out2(58,11);
	s_locks_lower_in(57,10) <= s_locks_lower_out(58,10);

		normal_cell_57_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,11),
			fetch              => s_fetch(57,11),
			data_in            => s_data_in(57,11),
			data_out           => s_data_out(57,11),
			out1               => s_out1(57,11),
			out2               => s_out2(57,11),
			lock_lower_row_out => s_locks_lower_out(57,11),
			lock_lower_row_in  => s_locks_lower_in(57,11),
			in1                => s_in1(57,11),
			in2                => s_in2(57,11),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(11)
		);
	s_in1(57,11)            <= s_out1(58,11);
	s_in2(57,11)            <= s_out2(58,12);
	s_locks_lower_in(57,11) <= s_locks_lower_out(58,11);

		normal_cell_57_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,12),
			fetch              => s_fetch(57,12),
			data_in            => s_data_in(57,12),
			data_out           => s_data_out(57,12),
			out1               => s_out1(57,12),
			out2               => s_out2(57,12),
			lock_lower_row_out => s_locks_lower_out(57,12),
			lock_lower_row_in  => s_locks_lower_in(57,12),
			in1                => s_in1(57,12),
			in2                => s_in2(57,12),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(12)
		);
	s_in1(57,12)            <= s_out1(58,12);
	s_in2(57,12)            <= s_out2(58,13);
	s_locks_lower_in(57,12) <= s_locks_lower_out(58,12);

		normal_cell_57_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,13),
			fetch              => s_fetch(57,13),
			data_in            => s_data_in(57,13),
			data_out           => s_data_out(57,13),
			out1               => s_out1(57,13),
			out2               => s_out2(57,13),
			lock_lower_row_out => s_locks_lower_out(57,13),
			lock_lower_row_in  => s_locks_lower_in(57,13),
			in1                => s_in1(57,13),
			in2                => s_in2(57,13),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(13)
		);
	s_in1(57,13)            <= s_out1(58,13);
	s_in2(57,13)            <= s_out2(58,14);
	s_locks_lower_in(57,13) <= s_locks_lower_out(58,13);

		normal_cell_57_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,14),
			fetch              => s_fetch(57,14),
			data_in            => s_data_in(57,14),
			data_out           => s_data_out(57,14),
			out1               => s_out1(57,14),
			out2               => s_out2(57,14),
			lock_lower_row_out => s_locks_lower_out(57,14),
			lock_lower_row_in  => s_locks_lower_in(57,14),
			in1                => s_in1(57,14),
			in2                => s_in2(57,14),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(14)
		);
	s_in1(57,14)            <= s_out1(58,14);
	s_in2(57,14)            <= s_out2(58,15);
	s_locks_lower_in(57,14) <= s_locks_lower_out(58,14);

		normal_cell_57_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,15),
			fetch              => s_fetch(57,15),
			data_in            => s_data_in(57,15),
			data_out           => s_data_out(57,15),
			out1               => s_out1(57,15),
			out2               => s_out2(57,15),
			lock_lower_row_out => s_locks_lower_out(57,15),
			lock_lower_row_in  => s_locks_lower_in(57,15),
			in1                => s_in1(57,15),
			in2                => s_in2(57,15),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(15)
		);
	s_in1(57,15)            <= s_out1(58,15);
	s_in2(57,15)            <= s_out2(58,16);
	s_locks_lower_in(57,15) <= s_locks_lower_out(58,15);

		normal_cell_57_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,16),
			fetch              => s_fetch(57,16),
			data_in            => s_data_in(57,16),
			data_out           => s_data_out(57,16),
			out1               => s_out1(57,16),
			out2               => s_out2(57,16),
			lock_lower_row_out => s_locks_lower_out(57,16),
			lock_lower_row_in  => s_locks_lower_in(57,16),
			in1                => s_in1(57,16),
			in2                => s_in2(57,16),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(16)
		);
	s_in1(57,16)            <= s_out1(58,16);
	s_in2(57,16)            <= s_out2(58,17);
	s_locks_lower_in(57,16) <= s_locks_lower_out(58,16);

		normal_cell_57_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,17),
			fetch              => s_fetch(57,17),
			data_in            => s_data_in(57,17),
			data_out           => s_data_out(57,17),
			out1               => s_out1(57,17),
			out2               => s_out2(57,17),
			lock_lower_row_out => s_locks_lower_out(57,17),
			lock_lower_row_in  => s_locks_lower_in(57,17),
			in1                => s_in1(57,17),
			in2                => s_in2(57,17),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(17)
		);
	s_in1(57,17)            <= s_out1(58,17);
	s_in2(57,17)            <= s_out2(58,18);
	s_locks_lower_in(57,17) <= s_locks_lower_out(58,17);

		normal_cell_57_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,18),
			fetch              => s_fetch(57,18),
			data_in            => s_data_in(57,18),
			data_out           => s_data_out(57,18),
			out1               => s_out1(57,18),
			out2               => s_out2(57,18),
			lock_lower_row_out => s_locks_lower_out(57,18),
			lock_lower_row_in  => s_locks_lower_in(57,18),
			in1                => s_in1(57,18),
			in2                => s_in2(57,18),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(18)
		);
	s_in1(57,18)            <= s_out1(58,18);
	s_in2(57,18)            <= s_out2(58,19);
	s_locks_lower_in(57,18) <= s_locks_lower_out(58,18);

		normal_cell_57_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,19),
			fetch              => s_fetch(57,19),
			data_in            => s_data_in(57,19),
			data_out           => s_data_out(57,19),
			out1               => s_out1(57,19),
			out2               => s_out2(57,19),
			lock_lower_row_out => s_locks_lower_out(57,19),
			lock_lower_row_in  => s_locks_lower_in(57,19),
			in1                => s_in1(57,19),
			in2                => s_in2(57,19),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(19)
		);
	s_in1(57,19)            <= s_out1(58,19);
	s_in2(57,19)            <= s_out2(58,20);
	s_locks_lower_in(57,19) <= s_locks_lower_out(58,19);

		normal_cell_57_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,20),
			fetch              => s_fetch(57,20),
			data_in            => s_data_in(57,20),
			data_out           => s_data_out(57,20),
			out1               => s_out1(57,20),
			out2               => s_out2(57,20),
			lock_lower_row_out => s_locks_lower_out(57,20),
			lock_lower_row_in  => s_locks_lower_in(57,20),
			in1                => s_in1(57,20),
			in2                => s_in2(57,20),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(20)
		);
	s_in1(57,20)            <= s_out1(58,20);
	s_in2(57,20)            <= s_out2(58,21);
	s_locks_lower_in(57,20) <= s_locks_lower_out(58,20);

		normal_cell_57_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,21),
			fetch              => s_fetch(57,21),
			data_in            => s_data_in(57,21),
			data_out           => s_data_out(57,21),
			out1               => s_out1(57,21),
			out2               => s_out2(57,21),
			lock_lower_row_out => s_locks_lower_out(57,21),
			lock_lower_row_in  => s_locks_lower_in(57,21),
			in1                => s_in1(57,21),
			in2                => s_in2(57,21),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(21)
		);
	s_in1(57,21)            <= s_out1(58,21);
	s_in2(57,21)            <= s_out2(58,22);
	s_locks_lower_in(57,21) <= s_locks_lower_out(58,21);

		normal_cell_57_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,22),
			fetch              => s_fetch(57,22),
			data_in            => s_data_in(57,22),
			data_out           => s_data_out(57,22),
			out1               => s_out1(57,22),
			out2               => s_out2(57,22),
			lock_lower_row_out => s_locks_lower_out(57,22),
			lock_lower_row_in  => s_locks_lower_in(57,22),
			in1                => s_in1(57,22),
			in2                => s_in2(57,22),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(22)
		);
	s_in1(57,22)            <= s_out1(58,22);
	s_in2(57,22)            <= s_out2(58,23);
	s_locks_lower_in(57,22) <= s_locks_lower_out(58,22);

		normal_cell_57_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,23),
			fetch              => s_fetch(57,23),
			data_in            => s_data_in(57,23),
			data_out           => s_data_out(57,23),
			out1               => s_out1(57,23),
			out2               => s_out2(57,23),
			lock_lower_row_out => s_locks_lower_out(57,23),
			lock_lower_row_in  => s_locks_lower_in(57,23),
			in1                => s_in1(57,23),
			in2                => s_in2(57,23),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(23)
		);
	s_in1(57,23)            <= s_out1(58,23);
	s_in2(57,23)            <= s_out2(58,24);
	s_locks_lower_in(57,23) <= s_locks_lower_out(58,23);

		normal_cell_57_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,24),
			fetch              => s_fetch(57,24),
			data_in            => s_data_in(57,24),
			data_out           => s_data_out(57,24),
			out1               => s_out1(57,24),
			out2               => s_out2(57,24),
			lock_lower_row_out => s_locks_lower_out(57,24),
			lock_lower_row_in  => s_locks_lower_in(57,24),
			in1                => s_in1(57,24),
			in2                => s_in2(57,24),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(24)
		);
	s_in1(57,24)            <= s_out1(58,24);
	s_in2(57,24)            <= s_out2(58,25);
	s_locks_lower_in(57,24) <= s_locks_lower_out(58,24);

		normal_cell_57_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,25),
			fetch              => s_fetch(57,25),
			data_in            => s_data_in(57,25),
			data_out           => s_data_out(57,25),
			out1               => s_out1(57,25),
			out2               => s_out2(57,25),
			lock_lower_row_out => s_locks_lower_out(57,25),
			lock_lower_row_in  => s_locks_lower_in(57,25),
			in1                => s_in1(57,25),
			in2                => s_in2(57,25),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(25)
		);
	s_in1(57,25)            <= s_out1(58,25);
	s_in2(57,25)            <= s_out2(58,26);
	s_locks_lower_in(57,25) <= s_locks_lower_out(58,25);

		normal_cell_57_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,26),
			fetch              => s_fetch(57,26),
			data_in            => s_data_in(57,26),
			data_out           => s_data_out(57,26),
			out1               => s_out1(57,26),
			out2               => s_out2(57,26),
			lock_lower_row_out => s_locks_lower_out(57,26),
			lock_lower_row_in  => s_locks_lower_in(57,26),
			in1                => s_in1(57,26),
			in2                => s_in2(57,26),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(26)
		);
	s_in1(57,26)            <= s_out1(58,26);
	s_in2(57,26)            <= s_out2(58,27);
	s_locks_lower_in(57,26) <= s_locks_lower_out(58,26);

		normal_cell_57_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,27),
			fetch              => s_fetch(57,27),
			data_in            => s_data_in(57,27),
			data_out           => s_data_out(57,27),
			out1               => s_out1(57,27),
			out2               => s_out2(57,27),
			lock_lower_row_out => s_locks_lower_out(57,27),
			lock_lower_row_in  => s_locks_lower_in(57,27),
			in1                => s_in1(57,27),
			in2                => s_in2(57,27),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(27)
		);
	s_in1(57,27)            <= s_out1(58,27);
	s_in2(57,27)            <= s_out2(58,28);
	s_locks_lower_in(57,27) <= s_locks_lower_out(58,27);

		normal_cell_57_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,28),
			fetch              => s_fetch(57,28),
			data_in            => s_data_in(57,28),
			data_out           => s_data_out(57,28),
			out1               => s_out1(57,28),
			out2               => s_out2(57,28),
			lock_lower_row_out => s_locks_lower_out(57,28),
			lock_lower_row_in  => s_locks_lower_in(57,28),
			in1                => s_in1(57,28),
			in2                => s_in2(57,28),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(28)
		);
	s_in1(57,28)            <= s_out1(58,28);
	s_in2(57,28)            <= s_out2(58,29);
	s_locks_lower_in(57,28) <= s_locks_lower_out(58,28);

		normal_cell_57_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,29),
			fetch              => s_fetch(57,29),
			data_in            => s_data_in(57,29),
			data_out           => s_data_out(57,29),
			out1               => s_out1(57,29),
			out2               => s_out2(57,29),
			lock_lower_row_out => s_locks_lower_out(57,29),
			lock_lower_row_in  => s_locks_lower_in(57,29),
			in1                => s_in1(57,29),
			in2                => s_in2(57,29),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(29)
		);
	s_in1(57,29)            <= s_out1(58,29);
	s_in2(57,29)            <= s_out2(58,30);
	s_locks_lower_in(57,29) <= s_locks_lower_out(58,29);

		normal_cell_57_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,30),
			fetch              => s_fetch(57,30),
			data_in            => s_data_in(57,30),
			data_out           => s_data_out(57,30),
			out1               => s_out1(57,30),
			out2               => s_out2(57,30),
			lock_lower_row_out => s_locks_lower_out(57,30),
			lock_lower_row_in  => s_locks_lower_in(57,30),
			in1                => s_in1(57,30),
			in2                => s_in2(57,30),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(30)
		);
	s_in1(57,30)            <= s_out1(58,30);
	s_in2(57,30)            <= s_out2(58,31);
	s_locks_lower_in(57,30) <= s_locks_lower_out(58,30);

		normal_cell_57_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,31),
			fetch              => s_fetch(57,31),
			data_in            => s_data_in(57,31),
			data_out           => s_data_out(57,31),
			out1               => s_out1(57,31),
			out2               => s_out2(57,31),
			lock_lower_row_out => s_locks_lower_out(57,31),
			lock_lower_row_in  => s_locks_lower_in(57,31),
			in1                => s_in1(57,31),
			in2                => s_in2(57,31),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(31)
		);
	s_in1(57,31)            <= s_out1(58,31);
	s_in2(57,31)            <= s_out2(58,32);
	s_locks_lower_in(57,31) <= s_locks_lower_out(58,31);

		normal_cell_57_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,32),
			fetch              => s_fetch(57,32),
			data_in            => s_data_in(57,32),
			data_out           => s_data_out(57,32),
			out1               => s_out1(57,32),
			out2               => s_out2(57,32),
			lock_lower_row_out => s_locks_lower_out(57,32),
			lock_lower_row_in  => s_locks_lower_in(57,32),
			in1                => s_in1(57,32),
			in2                => s_in2(57,32),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(32)
		);
	s_in1(57,32)            <= s_out1(58,32);
	s_in2(57,32)            <= s_out2(58,33);
	s_locks_lower_in(57,32) <= s_locks_lower_out(58,32);

		normal_cell_57_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,33),
			fetch              => s_fetch(57,33),
			data_in            => s_data_in(57,33),
			data_out           => s_data_out(57,33),
			out1               => s_out1(57,33),
			out2               => s_out2(57,33),
			lock_lower_row_out => s_locks_lower_out(57,33),
			lock_lower_row_in  => s_locks_lower_in(57,33),
			in1                => s_in1(57,33),
			in2                => s_in2(57,33),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(33)
		);
	s_in1(57,33)            <= s_out1(58,33);
	s_in2(57,33)            <= s_out2(58,34);
	s_locks_lower_in(57,33) <= s_locks_lower_out(58,33);

		normal_cell_57_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,34),
			fetch              => s_fetch(57,34),
			data_in            => s_data_in(57,34),
			data_out           => s_data_out(57,34),
			out1               => s_out1(57,34),
			out2               => s_out2(57,34),
			lock_lower_row_out => s_locks_lower_out(57,34),
			lock_lower_row_in  => s_locks_lower_in(57,34),
			in1                => s_in1(57,34),
			in2                => s_in2(57,34),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(34)
		);
	s_in1(57,34)            <= s_out1(58,34);
	s_in2(57,34)            <= s_out2(58,35);
	s_locks_lower_in(57,34) <= s_locks_lower_out(58,34);

		normal_cell_57_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,35),
			fetch              => s_fetch(57,35),
			data_in            => s_data_in(57,35),
			data_out           => s_data_out(57,35),
			out1               => s_out1(57,35),
			out2               => s_out2(57,35),
			lock_lower_row_out => s_locks_lower_out(57,35),
			lock_lower_row_in  => s_locks_lower_in(57,35),
			in1                => s_in1(57,35),
			in2                => s_in2(57,35),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(35)
		);
	s_in1(57,35)            <= s_out1(58,35);
	s_in2(57,35)            <= s_out2(58,36);
	s_locks_lower_in(57,35) <= s_locks_lower_out(58,35);

		normal_cell_57_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,36),
			fetch              => s_fetch(57,36),
			data_in            => s_data_in(57,36),
			data_out           => s_data_out(57,36),
			out1               => s_out1(57,36),
			out2               => s_out2(57,36),
			lock_lower_row_out => s_locks_lower_out(57,36),
			lock_lower_row_in  => s_locks_lower_in(57,36),
			in1                => s_in1(57,36),
			in2                => s_in2(57,36),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(36)
		);
	s_in1(57,36)            <= s_out1(58,36);
	s_in2(57,36)            <= s_out2(58,37);
	s_locks_lower_in(57,36) <= s_locks_lower_out(58,36);

		normal_cell_57_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,37),
			fetch              => s_fetch(57,37),
			data_in            => s_data_in(57,37),
			data_out           => s_data_out(57,37),
			out1               => s_out1(57,37),
			out2               => s_out2(57,37),
			lock_lower_row_out => s_locks_lower_out(57,37),
			lock_lower_row_in  => s_locks_lower_in(57,37),
			in1                => s_in1(57,37),
			in2                => s_in2(57,37),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(37)
		);
	s_in1(57,37)            <= s_out1(58,37);
	s_in2(57,37)            <= s_out2(58,38);
	s_locks_lower_in(57,37) <= s_locks_lower_out(58,37);

		normal_cell_57_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,38),
			fetch              => s_fetch(57,38),
			data_in            => s_data_in(57,38),
			data_out           => s_data_out(57,38),
			out1               => s_out1(57,38),
			out2               => s_out2(57,38),
			lock_lower_row_out => s_locks_lower_out(57,38),
			lock_lower_row_in  => s_locks_lower_in(57,38),
			in1                => s_in1(57,38),
			in2                => s_in2(57,38),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(38)
		);
	s_in1(57,38)            <= s_out1(58,38);
	s_in2(57,38)            <= s_out2(58,39);
	s_locks_lower_in(57,38) <= s_locks_lower_out(58,38);

		normal_cell_57_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,39),
			fetch              => s_fetch(57,39),
			data_in            => s_data_in(57,39),
			data_out           => s_data_out(57,39),
			out1               => s_out1(57,39),
			out2               => s_out2(57,39),
			lock_lower_row_out => s_locks_lower_out(57,39),
			lock_lower_row_in  => s_locks_lower_in(57,39),
			in1                => s_in1(57,39),
			in2                => s_in2(57,39),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(39)
		);
	s_in1(57,39)            <= s_out1(58,39);
	s_in2(57,39)            <= s_out2(58,40);
	s_locks_lower_in(57,39) <= s_locks_lower_out(58,39);

		normal_cell_57_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,40),
			fetch              => s_fetch(57,40),
			data_in            => s_data_in(57,40),
			data_out           => s_data_out(57,40),
			out1               => s_out1(57,40),
			out2               => s_out2(57,40),
			lock_lower_row_out => s_locks_lower_out(57,40),
			lock_lower_row_in  => s_locks_lower_in(57,40),
			in1                => s_in1(57,40),
			in2                => s_in2(57,40),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(40)
		);
	s_in1(57,40)            <= s_out1(58,40);
	s_in2(57,40)            <= s_out2(58,41);
	s_locks_lower_in(57,40) <= s_locks_lower_out(58,40);

		normal_cell_57_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,41),
			fetch              => s_fetch(57,41),
			data_in            => s_data_in(57,41),
			data_out           => s_data_out(57,41),
			out1               => s_out1(57,41),
			out2               => s_out2(57,41),
			lock_lower_row_out => s_locks_lower_out(57,41),
			lock_lower_row_in  => s_locks_lower_in(57,41),
			in1                => s_in1(57,41),
			in2                => s_in2(57,41),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(41)
		);
	s_in1(57,41)            <= s_out1(58,41);
	s_in2(57,41)            <= s_out2(58,42);
	s_locks_lower_in(57,41) <= s_locks_lower_out(58,41);

		normal_cell_57_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,42),
			fetch              => s_fetch(57,42),
			data_in            => s_data_in(57,42),
			data_out           => s_data_out(57,42),
			out1               => s_out1(57,42),
			out2               => s_out2(57,42),
			lock_lower_row_out => s_locks_lower_out(57,42),
			lock_lower_row_in  => s_locks_lower_in(57,42),
			in1                => s_in1(57,42),
			in2                => s_in2(57,42),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(42)
		);
	s_in1(57,42)            <= s_out1(58,42);
	s_in2(57,42)            <= s_out2(58,43);
	s_locks_lower_in(57,42) <= s_locks_lower_out(58,42);

		normal_cell_57_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,43),
			fetch              => s_fetch(57,43),
			data_in            => s_data_in(57,43),
			data_out           => s_data_out(57,43),
			out1               => s_out1(57,43),
			out2               => s_out2(57,43),
			lock_lower_row_out => s_locks_lower_out(57,43),
			lock_lower_row_in  => s_locks_lower_in(57,43),
			in1                => s_in1(57,43),
			in2                => s_in2(57,43),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(43)
		);
	s_in1(57,43)            <= s_out1(58,43);
	s_in2(57,43)            <= s_out2(58,44);
	s_locks_lower_in(57,43) <= s_locks_lower_out(58,43);

		normal_cell_57_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,44),
			fetch              => s_fetch(57,44),
			data_in            => s_data_in(57,44),
			data_out           => s_data_out(57,44),
			out1               => s_out1(57,44),
			out2               => s_out2(57,44),
			lock_lower_row_out => s_locks_lower_out(57,44),
			lock_lower_row_in  => s_locks_lower_in(57,44),
			in1                => s_in1(57,44),
			in2                => s_in2(57,44),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(44)
		);
	s_in1(57,44)            <= s_out1(58,44);
	s_in2(57,44)            <= s_out2(58,45);
	s_locks_lower_in(57,44) <= s_locks_lower_out(58,44);

		normal_cell_57_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,45),
			fetch              => s_fetch(57,45),
			data_in            => s_data_in(57,45),
			data_out           => s_data_out(57,45),
			out1               => s_out1(57,45),
			out2               => s_out2(57,45),
			lock_lower_row_out => s_locks_lower_out(57,45),
			lock_lower_row_in  => s_locks_lower_in(57,45),
			in1                => s_in1(57,45),
			in2                => s_in2(57,45),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(45)
		);
	s_in1(57,45)            <= s_out1(58,45);
	s_in2(57,45)            <= s_out2(58,46);
	s_locks_lower_in(57,45) <= s_locks_lower_out(58,45);

		normal_cell_57_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,46),
			fetch              => s_fetch(57,46),
			data_in            => s_data_in(57,46),
			data_out           => s_data_out(57,46),
			out1               => s_out1(57,46),
			out2               => s_out2(57,46),
			lock_lower_row_out => s_locks_lower_out(57,46),
			lock_lower_row_in  => s_locks_lower_in(57,46),
			in1                => s_in1(57,46),
			in2                => s_in2(57,46),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(46)
		);
	s_in1(57,46)            <= s_out1(58,46);
	s_in2(57,46)            <= s_out2(58,47);
	s_locks_lower_in(57,46) <= s_locks_lower_out(58,46);

		normal_cell_57_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,47),
			fetch              => s_fetch(57,47),
			data_in            => s_data_in(57,47),
			data_out           => s_data_out(57,47),
			out1               => s_out1(57,47),
			out2               => s_out2(57,47),
			lock_lower_row_out => s_locks_lower_out(57,47),
			lock_lower_row_in  => s_locks_lower_in(57,47),
			in1                => s_in1(57,47),
			in2                => s_in2(57,47),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(47)
		);
	s_in1(57,47)            <= s_out1(58,47);
	s_in2(57,47)            <= s_out2(58,48);
	s_locks_lower_in(57,47) <= s_locks_lower_out(58,47);

		normal_cell_57_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,48),
			fetch              => s_fetch(57,48),
			data_in            => s_data_in(57,48),
			data_out           => s_data_out(57,48),
			out1               => s_out1(57,48),
			out2               => s_out2(57,48),
			lock_lower_row_out => s_locks_lower_out(57,48),
			lock_lower_row_in  => s_locks_lower_in(57,48),
			in1                => s_in1(57,48),
			in2                => s_in2(57,48),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(48)
		);
	s_in1(57,48)            <= s_out1(58,48);
	s_in2(57,48)            <= s_out2(58,49);
	s_locks_lower_in(57,48) <= s_locks_lower_out(58,48);

		normal_cell_57_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,49),
			fetch              => s_fetch(57,49),
			data_in            => s_data_in(57,49),
			data_out           => s_data_out(57,49),
			out1               => s_out1(57,49),
			out2               => s_out2(57,49),
			lock_lower_row_out => s_locks_lower_out(57,49),
			lock_lower_row_in  => s_locks_lower_in(57,49),
			in1                => s_in1(57,49),
			in2                => s_in2(57,49),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(49)
		);
	s_in1(57,49)            <= s_out1(58,49);
	s_in2(57,49)            <= s_out2(58,50);
	s_locks_lower_in(57,49) <= s_locks_lower_out(58,49);

		normal_cell_57_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,50),
			fetch              => s_fetch(57,50),
			data_in            => s_data_in(57,50),
			data_out           => s_data_out(57,50),
			out1               => s_out1(57,50),
			out2               => s_out2(57,50),
			lock_lower_row_out => s_locks_lower_out(57,50),
			lock_lower_row_in  => s_locks_lower_in(57,50),
			in1                => s_in1(57,50),
			in2                => s_in2(57,50),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(50)
		);
	s_in1(57,50)            <= s_out1(58,50);
	s_in2(57,50)            <= s_out2(58,51);
	s_locks_lower_in(57,50) <= s_locks_lower_out(58,50);

		normal_cell_57_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,51),
			fetch              => s_fetch(57,51),
			data_in            => s_data_in(57,51),
			data_out           => s_data_out(57,51),
			out1               => s_out1(57,51),
			out2               => s_out2(57,51),
			lock_lower_row_out => s_locks_lower_out(57,51),
			lock_lower_row_in  => s_locks_lower_in(57,51),
			in1                => s_in1(57,51),
			in2                => s_in2(57,51),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(51)
		);
	s_in1(57,51)            <= s_out1(58,51);
	s_in2(57,51)            <= s_out2(58,52);
	s_locks_lower_in(57,51) <= s_locks_lower_out(58,51);

		normal_cell_57_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,52),
			fetch              => s_fetch(57,52),
			data_in            => s_data_in(57,52),
			data_out           => s_data_out(57,52),
			out1               => s_out1(57,52),
			out2               => s_out2(57,52),
			lock_lower_row_out => s_locks_lower_out(57,52),
			lock_lower_row_in  => s_locks_lower_in(57,52),
			in1                => s_in1(57,52),
			in2                => s_in2(57,52),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(52)
		);
	s_in1(57,52)            <= s_out1(58,52);
	s_in2(57,52)            <= s_out2(58,53);
	s_locks_lower_in(57,52) <= s_locks_lower_out(58,52);

		normal_cell_57_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,53),
			fetch              => s_fetch(57,53),
			data_in            => s_data_in(57,53),
			data_out           => s_data_out(57,53),
			out1               => s_out1(57,53),
			out2               => s_out2(57,53),
			lock_lower_row_out => s_locks_lower_out(57,53),
			lock_lower_row_in  => s_locks_lower_in(57,53),
			in1                => s_in1(57,53),
			in2                => s_in2(57,53),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(53)
		);
	s_in1(57,53)            <= s_out1(58,53);
	s_in2(57,53)            <= s_out2(58,54);
	s_locks_lower_in(57,53) <= s_locks_lower_out(58,53);

		normal_cell_57_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,54),
			fetch              => s_fetch(57,54),
			data_in            => s_data_in(57,54),
			data_out           => s_data_out(57,54),
			out1               => s_out1(57,54),
			out2               => s_out2(57,54),
			lock_lower_row_out => s_locks_lower_out(57,54),
			lock_lower_row_in  => s_locks_lower_in(57,54),
			in1                => s_in1(57,54),
			in2                => s_in2(57,54),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(54)
		);
	s_in1(57,54)            <= s_out1(58,54);
	s_in2(57,54)            <= s_out2(58,55);
	s_locks_lower_in(57,54) <= s_locks_lower_out(58,54);

		normal_cell_57_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,55),
			fetch              => s_fetch(57,55),
			data_in            => s_data_in(57,55),
			data_out           => s_data_out(57,55),
			out1               => s_out1(57,55),
			out2               => s_out2(57,55),
			lock_lower_row_out => s_locks_lower_out(57,55),
			lock_lower_row_in  => s_locks_lower_in(57,55),
			in1                => s_in1(57,55),
			in2                => s_in2(57,55),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(55)
		);
	s_in1(57,55)            <= s_out1(58,55);
	s_in2(57,55)            <= s_out2(58,56);
	s_locks_lower_in(57,55) <= s_locks_lower_out(58,55);

		normal_cell_57_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,56),
			fetch              => s_fetch(57,56),
			data_in            => s_data_in(57,56),
			data_out           => s_data_out(57,56),
			out1               => s_out1(57,56),
			out2               => s_out2(57,56),
			lock_lower_row_out => s_locks_lower_out(57,56),
			lock_lower_row_in  => s_locks_lower_in(57,56),
			in1                => s_in1(57,56),
			in2                => s_in2(57,56),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(56)
		);
	s_in1(57,56)            <= s_out1(58,56);
	s_in2(57,56)            <= s_out2(58,57);
	s_locks_lower_in(57,56) <= s_locks_lower_out(58,56);

		normal_cell_57_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,57),
			fetch              => s_fetch(57,57),
			data_in            => s_data_in(57,57),
			data_out           => s_data_out(57,57),
			out1               => s_out1(57,57),
			out2               => s_out2(57,57),
			lock_lower_row_out => s_locks_lower_out(57,57),
			lock_lower_row_in  => s_locks_lower_in(57,57),
			in1                => s_in1(57,57),
			in2                => s_in2(57,57),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(57)
		);
	s_in1(57,57)            <= s_out1(58,57);
	s_in2(57,57)            <= s_out2(58,58);
	s_locks_lower_in(57,57) <= s_locks_lower_out(58,57);

		normal_cell_57_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,58),
			fetch              => s_fetch(57,58),
			data_in            => s_data_in(57,58),
			data_out           => s_data_out(57,58),
			out1               => s_out1(57,58),
			out2               => s_out2(57,58),
			lock_lower_row_out => s_locks_lower_out(57,58),
			lock_lower_row_in  => s_locks_lower_in(57,58),
			in1                => s_in1(57,58),
			in2                => s_in2(57,58),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(58)
		);
	s_in1(57,58)            <= s_out1(58,58);
	s_in2(57,58)            <= s_out2(58,59);
	s_locks_lower_in(57,58) <= s_locks_lower_out(58,58);

		normal_cell_57_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,59),
			fetch              => s_fetch(57,59),
			data_in            => s_data_in(57,59),
			data_out           => s_data_out(57,59),
			out1               => s_out1(57,59),
			out2               => s_out2(57,59),
			lock_lower_row_out => s_locks_lower_out(57,59),
			lock_lower_row_in  => s_locks_lower_in(57,59),
			in1                => s_in1(57,59),
			in2                => s_in2(57,59),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(59)
		);
	s_in1(57,59)            <= s_out1(58,59);
	s_in2(57,59)            <= s_out2(58,60);
	s_locks_lower_in(57,59) <= s_locks_lower_out(58,59);

		last_col_cell_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(57,60),
			fetch              => s_fetch(57,60),
			data_in            => s_data_in(57,60),
			data_out           => s_data_out(57,60),
			out1               => s_out1(57,60),
			out2               => s_out2(57,60),
			lock_lower_row_out => s_locks_lower_out(57,60),
			lock_lower_row_in  => s_locks_lower_in(57,60),
			in1                => s_in1(57,60),
			in2                => (others => '0'),
			lock_row           => s_locks(57),
			piv_found          => s_piv_found,
			row_data           => s_row_data(57),
			col_data           => s_col_data(60)
		);
	s_in1(57,60)            <= s_out1(58,60);
	s_locks_lower_in(57,60) <= s_locks_lower_out(58,60);

		normal_cell_58_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,1),
			fetch              => s_fetch(58,1),
			data_in            => s_data_in(58,1),
			data_out           => s_data_out(58,1),
			out1               => s_out1(58,1),
			out2               => s_out2(58,1),
			lock_lower_row_out => s_locks_lower_out(58,1),
			lock_lower_row_in  => s_locks_lower_in(58,1),
			in1                => s_in1(58,1),
			in2                => s_in2(58,1),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(1)
		);
	s_in1(58,1)            <= s_out1(59,1);
	s_in2(58,1)            <= s_out2(59,2);
	s_locks_lower_in(58,1) <= s_locks_lower_out(59,1);

		normal_cell_58_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,2),
			fetch              => s_fetch(58,2),
			data_in            => s_data_in(58,2),
			data_out           => s_data_out(58,2),
			out1               => s_out1(58,2),
			out2               => s_out2(58,2),
			lock_lower_row_out => s_locks_lower_out(58,2),
			lock_lower_row_in  => s_locks_lower_in(58,2),
			in1                => s_in1(58,2),
			in2                => s_in2(58,2),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(2)
		);
	s_in1(58,2)            <= s_out1(59,2);
	s_in2(58,2)            <= s_out2(59,3);
	s_locks_lower_in(58,2) <= s_locks_lower_out(59,2);

		normal_cell_58_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,3),
			fetch              => s_fetch(58,3),
			data_in            => s_data_in(58,3),
			data_out           => s_data_out(58,3),
			out1               => s_out1(58,3),
			out2               => s_out2(58,3),
			lock_lower_row_out => s_locks_lower_out(58,3),
			lock_lower_row_in  => s_locks_lower_in(58,3),
			in1                => s_in1(58,3),
			in2                => s_in2(58,3),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(3)
		);
	s_in1(58,3)            <= s_out1(59,3);
	s_in2(58,3)            <= s_out2(59,4);
	s_locks_lower_in(58,3) <= s_locks_lower_out(59,3);

		normal_cell_58_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,4),
			fetch              => s_fetch(58,4),
			data_in            => s_data_in(58,4),
			data_out           => s_data_out(58,4),
			out1               => s_out1(58,4),
			out2               => s_out2(58,4),
			lock_lower_row_out => s_locks_lower_out(58,4),
			lock_lower_row_in  => s_locks_lower_in(58,4),
			in1                => s_in1(58,4),
			in2                => s_in2(58,4),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(4)
		);
	s_in1(58,4)            <= s_out1(59,4);
	s_in2(58,4)            <= s_out2(59,5);
	s_locks_lower_in(58,4) <= s_locks_lower_out(59,4);

		normal_cell_58_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,5),
			fetch              => s_fetch(58,5),
			data_in            => s_data_in(58,5),
			data_out           => s_data_out(58,5),
			out1               => s_out1(58,5),
			out2               => s_out2(58,5),
			lock_lower_row_out => s_locks_lower_out(58,5),
			lock_lower_row_in  => s_locks_lower_in(58,5),
			in1                => s_in1(58,5),
			in2                => s_in2(58,5),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(5)
		);
	s_in1(58,5)            <= s_out1(59,5);
	s_in2(58,5)            <= s_out2(59,6);
	s_locks_lower_in(58,5) <= s_locks_lower_out(59,5);

		normal_cell_58_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,6),
			fetch              => s_fetch(58,6),
			data_in            => s_data_in(58,6),
			data_out           => s_data_out(58,6),
			out1               => s_out1(58,6),
			out2               => s_out2(58,6),
			lock_lower_row_out => s_locks_lower_out(58,6),
			lock_lower_row_in  => s_locks_lower_in(58,6),
			in1                => s_in1(58,6),
			in2                => s_in2(58,6),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(6)
		);
	s_in1(58,6)            <= s_out1(59,6);
	s_in2(58,6)            <= s_out2(59,7);
	s_locks_lower_in(58,6) <= s_locks_lower_out(59,6);

		normal_cell_58_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,7),
			fetch              => s_fetch(58,7),
			data_in            => s_data_in(58,7),
			data_out           => s_data_out(58,7),
			out1               => s_out1(58,7),
			out2               => s_out2(58,7),
			lock_lower_row_out => s_locks_lower_out(58,7),
			lock_lower_row_in  => s_locks_lower_in(58,7),
			in1                => s_in1(58,7),
			in2                => s_in2(58,7),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(7)
		);
	s_in1(58,7)            <= s_out1(59,7);
	s_in2(58,7)            <= s_out2(59,8);
	s_locks_lower_in(58,7) <= s_locks_lower_out(59,7);

		normal_cell_58_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,8),
			fetch              => s_fetch(58,8),
			data_in            => s_data_in(58,8),
			data_out           => s_data_out(58,8),
			out1               => s_out1(58,8),
			out2               => s_out2(58,8),
			lock_lower_row_out => s_locks_lower_out(58,8),
			lock_lower_row_in  => s_locks_lower_in(58,8),
			in1                => s_in1(58,8),
			in2                => s_in2(58,8),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(8)
		);
	s_in1(58,8)            <= s_out1(59,8);
	s_in2(58,8)            <= s_out2(59,9);
	s_locks_lower_in(58,8) <= s_locks_lower_out(59,8);

		normal_cell_58_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,9),
			fetch              => s_fetch(58,9),
			data_in            => s_data_in(58,9),
			data_out           => s_data_out(58,9),
			out1               => s_out1(58,9),
			out2               => s_out2(58,9),
			lock_lower_row_out => s_locks_lower_out(58,9),
			lock_lower_row_in  => s_locks_lower_in(58,9),
			in1                => s_in1(58,9),
			in2                => s_in2(58,9),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(9)
		);
	s_in1(58,9)            <= s_out1(59,9);
	s_in2(58,9)            <= s_out2(59,10);
	s_locks_lower_in(58,9) <= s_locks_lower_out(59,9);

		normal_cell_58_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,10),
			fetch              => s_fetch(58,10),
			data_in            => s_data_in(58,10),
			data_out           => s_data_out(58,10),
			out1               => s_out1(58,10),
			out2               => s_out2(58,10),
			lock_lower_row_out => s_locks_lower_out(58,10),
			lock_lower_row_in  => s_locks_lower_in(58,10),
			in1                => s_in1(58,10),
			in2                => s_in2(58,10),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(10)
		);
	s_in1(58,10)            <= s_out1(59,10);
	s_in2(58,10)            <= s_out2(59,11);
	s_locks_lower_in(58,10) <= s_locks_lower_out(59,10);

		normal_cell_58_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,11),
			fetch              => s_fetch(58,11),
			data_in            => s_data_in(58,11),
			data_out           => s_data_out(58,11),
			out1               => s_out1(58,11),
			out2               => s_out2(58,11),
			lock_lower_row_out => s_locks_lower_out(58,11),
			lock_lower_row_in  => s_locks_lower_in(58,11),
			in1                => s_in1(58,11),
			in2                => s_in2(58,11),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(11)
		);
	s_in1(58,11)            <= s_out1(59,11);
	s_in2(58,11)            <= s_out2(59,12);
	s_locks_lower_in(58,11) <= s_locks_lower_out(59,11);

		normal_cell_58_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,12),
			fetch              => s_fetch(58,12),
			data_in            => s_data_in(58,12),
			data_out           => s_data_out(58,12),
			out1               => s_out1(58,12),
			out2               => s_out2(58,12),
			lock_lower_row_out => s_locks_lower_out(58,12),
			lock_lower_row_in  => s_locks_lower_in(58,12),
			in1                => s_in1(58,12),
			in2                => s_in2(58,12),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(12)
		);
	s_in1(58,12)            <= s_out1(59,12);
	s_in2(58,12)            <= s_out2(59,13);
	s_locks_lower_in(58,12) <= s_locks_lower_out(59,12);

		normal_cell_58_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,13),
			fetch              => s_fetch(58,13),
			data_in            => s_data_in(58,13),
			data_out           => s_data_out(58,13),
			out1               => s_out1(58,13),
			out2               => s_out2(58,13),
			lock_lower_row_out => s_locks_lower_out(58,13),
			lock_lower_row_in  => s_locks_lower_in(58,13),
			in1                => s_in1(58,13),
			in2                => s_in2(58,13),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(13)
		);
	s_in1(58,13)            <= s_out1(59,13);
	s_in2(58,13)            <= s_out2(59,14);
	s_locks_lower_in(58,13) <= s_locks_lower_out(59,13);

		normal_cell_58_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,14),
			fetch              => s_fetch(58,14),
			data_in            => s_data_in(58,14),
			data_out           => s_data_out(58,14),
			out1               => s_out1(58,14),
			out2               => s_out2(58,14),
			lock_lower_row_out => s_locks_lower_out(58,14),
			lock_lower_row_in  => s_locks_lower_in(58,14),
			in1                => s_in1(58,14),
			in2                => s_in2(58,14),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(14)
		);
	s_in1(58,14)            <= s_out1(59,14);
	s_in2(58,14)            <= s_out2(59,15);
	s_locks_lower_in(58,14) <= s_locks_lower_out(59,14);

		normal_cell_58_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,15),
			fetch              => s_fetch(58,15),
			data_in            => s_data_in(58,15),
			data_out           => s_data_out(58,15),
			out1               => s_out1(58,15),
			out2               => s_out2(58,15),
			lock_lower_row_out => s_locks_lower_out(58,15),
			lock_lower_row_in  => s_locks_lower_in(58,15),
			in1                => s_in1(58,15),
			in2                => s_in2(58,15),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(15)
		);
	s_in1(58,15)            <= s_out1(59,15);
	s_in2(58,15)            <= s_out2(59,16);
	s_locks_lower_in(58,15) <= s_locks_lower_out(59,15);

		normal_cell_58_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,16),
			fetch              => s_fetch(58,16),
			data_in            => s_data_in(58,16),
			data_out           => s_data_out(58,16),
			out1               => s_out1(58,16),
			out2               => s_out2(58,16),
			lock_lower_row_out => s_locks_lower_out(58,16),
			lock_lower_row_in  => s_locks_lower_in(58,16),
			in1                => s_in1(58,16),
			in2                => s_in2(58,16),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(16)
		);
	s_in1(58,16)            <= s_out1(59,16);
	s_in2(58,16)            <= s_out2(59,17);
	s_locks_lower_in(58,16) <= s_locks_lower_out(59,16);

		normal_cell_58_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,17),
			fetch              => s_fetch(58,17),
			data_in            => s_data_in(58,17),
			data_out           => s_data_out(58,17),
			out1               => s_out1(58,17),
			out2               => s_out2(58,17),
			lock_lower_row_out => s_locks_lower_out(58,17),
			lock_lower_row_in  => s_locks_lower_in(58,17),
			in1                => s_in1(58,17),
			in2                => s_in2(58,17),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(17)
		);
	s_in1(58,17)            <= s_out1(59,17);
	s_in2(58,17)            <= s_out2(59,18);
	s_locks_lower_in(58,17) <= s_locks_lower_out(59,17);

		normal_cell_58_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,18),
			fetch              => s_fetch(58,18),
			data_in            => s_data_in(58,18),
			data_out           => s_data_out(58,18),
			out1               => s_out1(58,18),
			out2               => s_out2(58,18),
			lock_lower_row_out => s_locks_lower_out(58,18),
			lock_lower_row_in  => s_locks_lower_in(58,18),
			in1                => s_in1(58,18),
			in2                => s_in2(58,18),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(18)
		);
	s_in1(58,18)            <= s_out1(59,18);
	s_in2(58,18)            <= s_out2(59,19);
	s_locks_lower_in(58,18) <= s_locks_lower_out(59,18);

		normal_cell_58_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,19),
			fetch              => s_fetch(58,19),
			data_in            => s_data_in(58,19),
			data_out           => s_data_out(58,19),
			out1               => s_out1(58,19),
			out2               => s_out2(58,19),
			lock_lower_row_out => s_locks_lower_out(58,19),
			lock_lower_row_in  => s_locks_lower_in(58,19),
			in1                => s_in1(58,19),
			in2                => s_in2(58,19),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(19)
		);
	s_in1(58,19)            <= s_out1(59,19);
	s_in2(58,19)            <= s_out2(59,20);
	s_locks_lower_in(58,19) <= s_locks_lower_out(59,19);

		normal_cell_58_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,20),
			fetch              => s_fetch(58,20),
			data_in            => s_data_in(58,20),
			data_out           => s_data_out(58,20),
			out1               => s_out1(58,20),
			out2               => s_out2(58,20),
			lock_lower_row_out => s_locks_lower_out(58,20),
			lock_lower_row_in  => s_locks_lower_in(58,20),
			in1                => s_in1(58,20),
			in2                => s_in2(58,20),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(20)
		);
	s_in1(58,20)            <= s_out1(59,20);
	s_in2(58,20)            <= s_out2(59,21);
	s_locks_lower_in(58,20) <= s_locks_lower_out(59,20);

		normal_cell_58_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,21),
			fetch              => s_fetch(58,21),
			data_in            => s_data_in(58,21),
			data_out           => s_data_out(58,21),
			out1               => s_out1(58,21),
			out2               => s_out2(58,21),
			lock_lower_row_out => s_locks_lower_out(58,21),
			lock_lower_row_in  => s_locks_lower_in(58,21),
			in1                => s_in1(58,21),
			in2                => s_in2(58,21),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(21)
		);
	s_in1(58,21)            <= s_out1(59,21);
	s_in2(58,21)            <= s_out2(59,22);
	s_locks_lower_in(58,21) <= s_locks_lower_out(59,21);

		normal_cell_58_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,22),
			fetch              => s_fetch(58,22),
			data_in            => s_data_in(58,22),
			data_out           => s_data_out(58,22),
			out1               => s_out1(58,22),
			out2               => s_out2(58,22),
			lock_lower_row_out => s_locks_lower_out(58,22),
			lock_lower_row_in  => s_locks_lower_in(58,22),
			in1                => s_in1(58,22),
			in2                => s_in2(58,22),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(22)
		);
	s_in1(58,22)            <= s_out1(59,22);
	s_in2(58,22)            <= s_out2(59,23);
	s_locks_lower_in(58,22) <= s_locks_lower_out(59,22);

		normal_cell_58_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,23),
			fetch              => s_fetch(58,23),
			data_in            => s_data_in(58,23),
			data_out           => s_data_out(58,23),
			out1               => s_out1(58,23),
			out2               => s_out2(58,23),
			lock_lower_row_out => s_locks_lower_out(58,23),
			lock_lower_row_in  => s_locks_lower_in(58,23),
			in1                => s_in1(58,23),
			in2                => s_in2(58,23),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(23)
		);
	s_in1(58,23)            <= s_out1(59,23);
	s_in2(58,23)            <= s_out2(59,24);
	s_locks_lower_in(58,23) <= s_locks_lower_out(59,23);

		normal_cell_58_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,24),
			fetch              => s_fetch(58,24),
			data_in            => s_data_in(58,24),
			data_out           => s_data_out(58,24),
			out1               => s_out1(58,24),
			out2               => s_out2(58,24),
			lock_lower_row_out => s_locks_lower_out(58,24),
			lock_lower_row_in  => s_locks_lower_in(58,24),
			in1                => s_in1(58,24),
			in2                => s_in2(58,24),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(24)
		);
	s_in1(58,24)            <= s_out1(59,24);
	s_in2(58,24)            <= s_out2(59,25);
	s_locks_lower_in(58,24) <= s_locks_lower_out(59,24);

		normal_cell_58_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,25),
			fetch              => s_fetch(58,25),
			data_in            => s_data_in(58,25),
			data_out           => s_data_out(58,25),
			out1               => s_out1(58,25),
			out2               => s_out2(58,25),
			lock_lower_row_out => s_locks_lower_out(58,25),
			lock_lower_row_in  => s_locks_lower_in(58,25),
			in1                => s_in1(58,25),
			in2                => s_in2(58,25),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(25)
		);
	s_in1(58,25)            <= s_out1(59,25);
	s_in2(58,25)            <= s_out2(59,26);
	s_locks_lower_in(58,25) <= s_locks_lower_out(59,25);

		normal_cell_58_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,26),
			fetch              => s_fetch(58,26),
			data_in            => s_data_in(58,26),
			data_out           => s_data_out(58,26),
			out1               => s_out1(58,26),
			out2               => s_out2(58,26),
			lock_lower_row_out => s_locks_lower_out(58,26),
			lock_lower_row_in  => s_locks_lower_in(58,26),
			in1                => s_in1(58,26),
			in2                => s_in2(58,26),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(26)
		);
	s_in1(58,26)            <= s_out1(59,26);
	s_in2(58,26)            <= s_out2(59,27);
	s_locks_lower_in(58,26) <= s_locks_lower_out(59,26);

		normal_cell_58_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,27),
			fetch              => s_fetch(58,27),
			data_in            => s_data_in(58,27),
			data_out           => s_data_out(58,27),
			out1               => s_out1(58,27),
			out2               => s_out2(58,27),
			lock_lower_row_out => s_locks_lower_out(58,27),
			lock_lower_row_in  => s_locks_lower_in(58,27),
			in1                => s_in1(58,27),
			in2                => s_in2(58,27),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(27)
		);
	s_in1(58,27)            <= s_out1(59,27);
	s_in2(58,27)            <= s_out2(59,28);
	s_locks_lower_in(58,27) <= s_locks_lower_out(59,27);

		normal_cell_58_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,28),
			fetch              => s_fetch(58,28),
			data_in            => s_data_in(58,28),
			data_out           => s_data_out(58,28),
			out1               => s_out1(58,28),
			out2               => s_out2(58,28),
			lock_lower_row_out => s_locks_lower_out(58,28),
			lock_lower_row_in  => s_locks_lower_in(58,28),
			in1                => s_in1(58,28),
			in2                => s_in2(58,28),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(28)
		);
	s_in1(58,28)            <= s_out1(59,28);
	s_in2(58,28)            <= s_out2(59,29);
	s_locks_lower_in(58,28) <= s_locks_lower_out(59,28);

		normal_cell_58_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,29),
			fetch              => s_fetch(58,29),
			data_in            => s_data_in(58,29),
			data_out           => s_data_out(58,29),
			out1               => s_out1(58,29),
			out2               => s_out2(58,29),
			lock_lower_row_out => s_locks_lower_out(58,29),
			lock_lower_row_in  => s_locks_lower_in(58,29),
			in1                => s_in1(58,29),
			in2                => s_in2(58,29),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(29)
		);
	s_in1(58,29)            <= s_out1(59,29);
	s_in2(58,29)            <= s_out2(59,30);
	s_locks_lower_in(58,29) <= s_locks_lower_out(59,29);

		normal_cell_58_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,30),
			fetch              => s_fetch(58,30),
			data_in            => s_data_in(58,30),
			data_out           => s_data_out(58,30),
			out1               => s_out1(58,30),
			out2               => s_out2(58,30),
			lock_lower_row_out => s_locks_lower_out(58,30),
			lock_lower_row_in  => s_locks_lower_in(58,30),
			in1                => s_in1(58,30),
			in2                => s_in2(58,30),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(30)
		);
	s_in1(58,30)            <= s_out1(59,30);
	s_in2(58,30)            <= s_out2(59,31);
	s_locks_lower_in(58,30) <= s_locks_lower_out(59,30);

		normal_cell_58_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,31),
			fetch              => s_fetch(58,31),
			data_in            => s_data_in(58,31),
			data_out           => s_data_out(58,31),
			out1               => s_out1(58,31),
			out2               => s_out2(58,31),
			lock_lower_row_out => s_locks_lower_out(58,31),
			lock_lower_row_in  => s_locks_lower_in(58,31),
			in1                => s_in1(58,31),
			in2                => s_in2(58,31),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(31)
		);
	s_in1(58,31)            <= s_out1(59,31);
	s_in2(58,31)            <= s_out2(59,32);
	s_locks_lower_in(58,31) <= s_locks_lower_out(59,31);

		normal_cell_58_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,32),
			fetch              => s_fetch(58,32),
			data_in            => s_data_in(58,32),
			data_out           => s_data_out(58,32),
			out1               => s_out1(58,32),
			out2               => s_out2(58,32),
			lock_lower_row_out => s_locks_lower_out(58,32),
			lock_lower_row_in  => s_locks_lower_in(58,32),
			in1                => s_in1(58,32),
			in2                => s_in2(58,32),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(32)
		);
	s_in1(58,32)            <= s_out1(59,32);
	s_in2(58,32)            <= s_out2(59,33);
	s_locks_lower_in(58,32) <= s_locks_lower_out(59,32);

		normal_cell_58_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,33),
			fetch              => s_fetch(58,33),
			data_in            => s_data_in(58,33),
			data_out           => s_data_out(58,33),
			out1               => s_out1(58,33),
			out2               => s_out2(58,33),
			lock_lower_row_out => s_locks_lower_out(58,33),
			lock_lower_row_in  => s_locks_lower_in(58,33),
			in1                => s_in1(58,33),
			in2                => s_in2(58,33),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(33)
		);
	s_in1(58,33)            <= s_out1(59,33);
	s_in2(58,33)            <= s_out2(59,34);
	s_locks_lower_in(58,33) <= s_locks_lower_out(59,33);

		normal_cell_58_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,34),
			fetch              => s_fetch(58,34),
			data_in            => s_data_in(58,34),
			data_out           => s_data_out(58,34),
			out1               => s_out1(58,34),
			out2               => s_out2(58,34),
			lock_lower_row_out => s_locks_lower_out(58,34),
			lock_lower_row_in  => s_locks_lower_in(58,34),
			in1                => s_in1(58,34),
			in2                => s_in2(58,34),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(34)
		);
	s_in1(58,34)            <= s_out1(59,34);
	s_in2(58,34)            <= s_out2(59,35);
	s_locks_lower_in(58,34) <= s_locks_lower_out(59,34);

		normal_cell_58_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,35),
			fetch              => s_fetch(58,35),
			data_in            => s_data_in(58,35),
			data_out           => s_data_out(58,35),
			out1               => s_out1(58,35),
			out2               => s_out2(58,35),
			lock_lower_row_out => s_locks_lower_out(58,35),
			lock_lower_row_in  => s_locks_lower_in(58,35),
			in1                => s_in1(58,35),
			in2                => s_in2(58,35),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(35)
		);
	s_in1(58,35)            <= s_out1(59,35);
	s_in2(58,35)            <= s_out2(59,36);
	s_locks_lower_in(58,35) <= s_locks_lower_out(59,35);

		normal_cell_58_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,36),
			fetch              => s_fetch(58,36),
			data_in            => s_data_in(58,36),
			data_out           => s_data_out(58,36),
			out1               => s_out1(58,36),
			out2               => s_out2(58,36),
			lock_lower_row_out => s_locks_lower_out(58,36),
			lock_lower_row_in  => s_locks_lower_in(58,36),
			in1                => s_in1(58,36),
			in2                => s_in2(58,36),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(36)
		);
	s_in1(58,36)            <= s_out1(59,36);
	s_in2(58,36)            <= s_out2(59,37);
	s_locks_lower_in(58,36) <= s_locks_lower_out(59,36);

		normal_cell_58_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,37),
			fetch              => s_fetch(58,37),
			data_in            => s_data_in(58,37),
			data_out           => s_data_out(58,37),
			out1               => s_out1(58,37),
			out2               => s_out2(58,37),
			lock_lower_row_out => s_locks_lower_out(58,37),
			lock_lower_row_in  => s_locks_lower_in(58,37),
			in1                => s_in1(58,37),
			in2                => s_in2(58,37),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(37)
		);
	s_in1(58,37)            <= s_out1(59,37);
	s_in2(58,37)            <= s_out2(59,38);
	s_locks_lower_in(58,37) <= s_locks_lower_out(59,37);

		normal_cell_58_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,38),
			fetch              => s_fetch(58,38),
			data_in            => s_data_in(58,38),
			data_out           => s_data_out(58,38),
			out1               => s_out1(58,38),
			out2               => s_out2(58,38),
			lock_lower_row_out => s_locks_lower_out(58,38),
			lock_lower_row_in  => s_locks_lower_in(58,38),
			in1                => s_in1(58,38),
			in2                => s_in2(58,38),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(38)
		);
	s_in1(58,38)            <= s_out1(59,38);
	s_in2(58,38)            <= s_out2(59,39);
	s_locks_lower_in(58,38) <= s_locks_lower_out(59,38);

		normal_cell_58_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,39),
			fetch              => s_fetch(58,39),
			data_in            => s_data_in(58,39),
			data_out           => s_data_out(58,39),
			out1               => s_out1(58,39),
			out2               => s_out2(58,39),
			lock_lower_row_out => s_locks_lower_out(58,39),
			lock_lower_row_in  => s_locks_lower_in(58,39),
			in1                => s_in1(58,39),
			in2                => s_in2(58,39),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(39)
		);
	s_in1(58,39)            <= s_out1(59,39);
	s_in2(58,39)            <= s_out2(59,40);
	s_locks_lower_in(58,39) <= s_locks_lower_out(59,39);

		normal_cell_58_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,40),
			fetch              => s_fetch(58,40),
			data_in            => s_data_in(58,40),
			data_out           => s_data_out(58,40),
			out1               => s_out1(58,40),
			out2               => s_out2(58,40),
			lock_lower_row_out => s_locks_lower_out(58,40),
			lock_lower_row_in  => s_locks_lower_in(58,40),
			in1                => s_in1(58,40),
			in2                => s_in2(58,40),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(40)
		);
	s_in1(58,40)            <= s_out1(59,40);
	s_in2(58,40)            <= s_out2(59,41);
	s_locks_lower_in(58,40) <= s_locks_lower_out(59,40);

		normal_cell_58_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,41),
			fetch              => s_fetch(58,41),
			data_in            => s_data_in(58,41),
			data_out           => s_data_out(58,41),
			out1               => s_out1(58,41),
			out2               => s_out2(58,41),
			lock_lower_row_out => s_locks_lower_out(58,41),
			lock_lower_row_in  => s_locks_lower_in(58,41),
			in1                => s_in1(58,41),
			in2                => s_in2(58,41),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(41)
		);
	s_in1(58,41)            <= s_out1(59,41);
	s_in2(58,41)            <= s_out2(59,42);
	s_locks_lower_in(58,41) <= s_locks_lower_out(59,41);

		normal_cell_58_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,42),
			fetch              => s_fetch(58,42),
			data_in            => s_data_in(58,42),
			data_out           => s_data_out(58,42),
			out1               => s_out1(58,42),
			out2               => s_out2(58,42),
			lock_lower_row_out => s_locks_lower_out(58,42),
			lock_lower_row_in  => s_locks_lower_in(58,42),
			in1                => s_in1(58,42),
			in2                => s_in2(58,42),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(42)
		);
	s_in1(58,42)            <= s_out1(59,42);
	s_in2(58,42)            <= s_out2(59,43);
	s_locks_lower_in(58,42) <= s_locks_lower_out(59,42);

		normal_cell_58_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,43),
			fetch              => s_fetch(58,43),
			data_in            => s_data_in(58,43),
			data_out           => s_data_out(58,43),
			out1               => s_out1(58,43),
			out2               => s_out2(58,43),
			lock_lower_row_out => s_locks_lower_out(58,43),
			lock_lower_row_in  => s_locks_lower_in(58,43),
			in1                => s_in1(58,43),
			in2                => s_in2(58,43),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(43)
		);
	s_in1(58,43)            <= s_out1(59,43);
	s_in2(58,43)            <= s_out2(59,44);
	s_locks_lower_in(58,43) <= s_locks_lower_out(59,43);

		normal_cell_58_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,44),
			fetch              => s_fetch(58,44),
			data_in            => s_data_in(58,44),
			data_out           => s_data_out(58,44),
			out1               => s_out1(58,44),
			out2               => s_out2(58,44),
			lock_lower_row_out => s_locks_lower_out(58,44),
			lock_lower_row_in  => s_locks_lower_in(58,44),
			in1                => s_in1(58,44),
			in2                => s_in2(58,44),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(44)
		);
	s_in1(58,44)            <= s_out1(59,44);
	s_in2(58,44)            <= s_out2(59,45);
	s_locks_lower_in(58,44) <= s_locks_lower_out(59,44);

		normal_cell_58_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,45),
			fetch              => s_fetch(58,45),
			data_in            => s_data_in(58,45),
			data_out           => s_data_out(58,45),
			out1               => s_out1(58,45),
			out2               => s_out2(58,45),
			lock_lower_row_out => s_locks_lower_out(58,45),
			lock_lower_row_in  => s_locks_lower_in(58,45),
			in1                => s_in1(58,45),
			in2                => s_in2(58,45),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(45)
		);
	s_in1(58,45)            <= s_out1(59,45);
	s_in2(58,45)            <= s_out2(59,46);
	s_locks_lower_in(58,45) <= s_locks_lower_out(59,45);

		normal_cell_58_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,46),
			fetch              => s_fetch(58,46),
			data_in            => s_data_in(58,46),
			data_out           => s_data_out(58,46),
			out1               => s_out1(58,46),
			out2               => s_out2(58,46),
			lock_lower_row_out => s_locks_lower_out(58,46),
			lock_lower_row_in  => s_locks_lower_in(58,46),
			in1                => s_in1(58,46),
			in2                => s_in2(58,46),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(46)
		);
	s_in1(58,46)            <= s_out1(59,46);
	s_in2(58,46)            <= s_out2(59,47);
	s_locks_lower_in(58,46) <= s_locks_lower_out(59,46);

		normal_cell_58_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,47),
			fetch              => s_fetch(58,47),
			data_in            => s_data_in(58,47),
			data_out           => s_data_out(58,47),
			out1               => s_out1(58,47),
			out2               => s_out2(58,47),
			lock_lower_row_out => s_locks_lower_out(58,47),
			lock_lower_row_in  => s_locks_lower_in(58,47),
			in1                => s_in1(58,47),
			in2                => s_in2(58,47),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(47)
		);
	s_in1(58,47)            <= s_out1(59,47);
	s_in2(58,47)            <= s_out2(59,48);
	s_locks_lower_in(58,47) <= s_locks_lower_out(59,47);

		normal_cell_58_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,48),
			fetch              => s_fetch(58,48),
			data_in            => s_data_in(58,48),
			data_out           => s_data_out(58,48),
			out1               => s_out1(58,48),
			out2               => s_out2(58,48),
			lock_lower_row_out => s_locks_lower_out(58,48),
			lock_lower_row_in  => s_locks_lower_in(58,48),
			in1                => s_in1(58,48),
			in2                => s_in2(58,48),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(48)
		);
	s_in1(58,48)            <= s_out1(59,48);
	s_in2(58,48)            <= s_out2(59,49);
	s_locks_lower_in(58,48) <= s_locks_lower_out(59,48);

		normal_cell_58_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,49),
			fetch              => s_fetch(58,49),
			data_in            => s_data_in(58,49),
			data_out           => s_data_out(58,49),
			out1               => s_out1(58,49),
			out2               => s_out2(58,49),
			lock_lower_row_out => s_locks_lower_out(58,49),
			lock_lower_row_in  => s_locks_lower_in(58,49),
			in1                => s_in1(58,49),
			in2                => s_in2(58,49),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(49)
		);
	s_in1(58,49)            <= s_out1(59,49);
	s_in2(58,49)            <= s_out2(59,50);
	s_locks_lower_in(58,49) <= s_locks_lower_out(59,49);

		normal_cell_58_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,50),
			fetch              => s_fetch(58,50),
			data_in            => s_data_in(58,50),
			data_out           => s_data_out(58,50),
			out1               => s_out1(58,50),
			out2               => s_out2(58,50),
			lock_lower_row_out => s_locks_lower_out(58,50),
			lock_lower_row_in  => s_locks_lower_in(58,50),
			in1                => s_in1(58,50),
			in2                => s_in2(58,50),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(50)
		);
	s_in1(58,50)            <= s_out1(59,50);
	s_in2(58,50)            <= s_out2(59,51);
	s_locks_lower_in(58,50) <= s_locks_lower_out(59,50);

		normal_cell_58_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,51),
			fetch              => s_fetch(58,51),
			data_in            => s_data_in(58,51),
			data_out           => s_data_out(58,51),
			out1               => s_out1(58,51),
			out2               => s_out2(58,51),
			lock_lower_row_out => s_locks_lower_out(58,51),
			lock_lower_row_in  => s_locks_lower_in(58,51),
			in1                => s_in1(58,51),
			in2                => s_in2(58,51),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(51)
		);
	s_in1(58,51)            <= s_out1(59,51);
	s_in2(58,51)            <= s_out2(59,52);
	s_locks_lower_in(58,51) <= s_locks_lower_out(59,51);

		normal_cell_58_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,52),
			fetch              => s_fetch(58,52),
			data_in            => s_data_in(58,52),
			data_out           => s_data_out(58,52),
			out1               => s_out1(58,52),
			out2               => s_out2(58,52),
			lock_lower_row_out => s_locks_lower_out(58,52),
			lock_lower_row_in  => s_locks_lower_in(58,52),
			in1                => s_in1(58,52),
			in2                => s_in2(58,52),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(52)
		);
	s_in1(58,52)            <= s_out1(59,52);
	s_in2(58,52)            <= s_out2(59,53);
	s_locks_lower_in(58,52) <= s_locks_lower_out(59,52);

		normal_cell_58_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,53),
			fetch              => s_fetch(58,53),
			data_in            => s_data_in(58,53),
			data_out           => s_data_out(58,53),
			out1               => s_out1(58,53),
			out2               => s_out2(58,53),
			lock_lower_row_out => s_locks_lower_out(58,53),
			lock_lower_row_in  => s_locks_lower_in(58,53),
			in1                => s_in1(58,53),
			in2                => s_in2(58,53),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(53)
		);
	s_in1(58,53)            <= s_out1(59,53);
	s_in2(58,53)            <= s_out2(59,54);
	s_locks_lower_in(58,53) <= s_locks_lower_out(59,53);

		normal_cell_58_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,54),
			fetch              => s_fetch(58,54),
			data_in            => s_data_in(58,54),
			data_out           => s_data_out(58,54),
			out1               => s_out1(58,54),
			out2               => s_out2(58,54),
			lock_lower_row_out => s_locks_lower_out(58,54),
			lock_lower_row_in  => s_locks_lower_in(58,54),
			in1                => s_in1(58,54),
			in2                => s_in2(58,54),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(54)
		);
	s_in1(58,54)            <= s_out1(59,54);
	s_in2(58,54)            <= s_out2(59,55);
	s_locks_lower_in(58,54) <= s_locks_lower_out(59,54);

		normal_cell_58_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,55),
			fetch              => s_fetch(58,55),
			data_in            => s_data_in(58,55),
			data_out           => s_data_out(58,55),
			out1               => s_out1(58,55),
			out2               => s_out2(58,55),
			lock_lower_row_out => s_locks_lower_out(58,55),
			lock_lower_row_in  => s_locks_lower_in(58,55),
			in1                => s_in1(58,55),
			in2                => s_in2(58,55),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(55)
		);
	s_in1(58,55)            <= s_out1(59,55);
	s_in2(58,55)            <= s_out2(59,56);
	s_locks_lower_in(58,55) <= s_locks_lower_out(59,55);

		normal_cell_58_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,56),
			fetch              => s_fetch(58,56),
			data_in            => s_data_in(58,56),
			data_out           => s_data_out(58,56),
			out1               => s_out1(58,56),
			out2               => s_out2(58,56),
			lock_lower_row_out => s_locks_lower_out(58,56),
			lock_lower_row_in  => s_locks_lower_in(58,56),
			in1                => s_in1(58,56),
			in2                => s_in2(58,56),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(56)
		);
	s_in1(58,56)            <= s_out1(59,56);
	s_in2(58,56)            <= s_out2(59,57);
	s_locks_lower_in(58,56) <= s_locks_lower_out(59,56);

		normal_cell_58_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,57),
			fetch              => s_fetch(58,57),
			data_in            => s_data_in(58,57),
			data_out           => s_data_out(58,57),
			out1               => s_out1(58,57),
			out2               => s_out2(58,57),
			lock_lower_row_out => s_locks_lower_out(58,57),
			lock_lower_row_in  => s_locks_lower_in(58,57),
			in1                => s_in1(58,57),
			in2                => s_in2(58,57),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(57)
		);
	s_in1(58,57)            <= s_out1(59,57);
	s_in2(58,57)            <= s_out2(59,58);
	s_locks_lower_in(58,57) <= s_locks_lower_out(59,57);

		normal_cell_58_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,58),
			fetch              => s_fetch(58,58),
			data_in            => s_data_in(58,58),
			data_out           => s_data_out(58,58),
			out1               => s_out1(58,58),
			out2               => s_out2(58,58),
			lock_lower_row_out => s_locks_lower_out(58,58),
			lock_lower_row_in  => s_locks_lower_in(58,58),
			in1                => s_in1(58,58),
			in2                => s_in2(58,58),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(58)
		);
	s_in1(58,58)            <= s_out1(59,58);
	s_in2(58,58)            <= s_out2(59,59);
	s_locks_lower_in(58,58) <= s_locks_lower_out(59,58);

		normal_cell_58_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,59),
			fetch              => s_fetch(58,59),
			data_in            => s_data_in(58,59),
			data_out           => s_data_out(58,59),
			out1               => s_out1(58,59),
			out2               => s_out2(58,59),
			lock_lower_row_out => s_locks_lower_out(58,59),
			lock_lower_row_in  => s_locks_lower_in(58,59),
			in1                => s_in1(58,59),
			in2                => s_in2(58,59),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(59)
		);
	s_in1(58,59)            <= s_out1(59,59);
	s_in2(58,59)            <= s_out2(59,60);
	s_locks_lower_in(58,59) <= s_locks_lower_out(59,59);

		last_col_cell_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(58,60),
			fetch              => s_fetch(58,60),
			data_in            => s_data_in(58,60),
			data_out           => s_data_out(58,60),
			out1               => s_out1(58,60),
			out2               => s_out2(58,60),
			lock_lower_row_out => s_locks_lower_out(58,60),
			lock_lower_row_in  => s_locks_lower_in(58,60),
			in1                => s_in1(58,60),
			in2                => (others => '0'),
			lock_row           => s_locks(58),
			piv_found          => s_piv_found,
			row_data           => s_row_data(58),
			col_data           => s_col_data(60)
		);
	s_in1(58,60)            <= s_out1(59,60);
	s_locks_lower_in(58,60) <= s_locks_lower_out(59,60);

		last_row_cell_1 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,1),
			fetch              => s_fetch(59,1),
			data_in            => s_data_in(59,1),
			data_out           => s_data_out(59,1),
			out1               => s_out1(59,1),
			out2               => s_out2(59,1),
			lock_lower_row_out => s_locks_lower_out(59,1),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,1),
			in2                => s_in2(59,1),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(1)
		);
	s_in1(59,1) <= s_out1(0,1);
	s_in2(59,1) <= s_out2(0,2);

		last_row_cell_2 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,2),
			fetch              => s_fetch(59,2),
			data_in            => s_data_in(59,2),
			data_out           => s_data_out(59,2),
			out1               => s_out1(59,2),
			out2               => s_out2(59,2),
			lock_lower_row_out => s_locks_lower_out(59,2),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,2),
			in2                => s_in2(59,2),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(2)
		);
	s_in1(59,2) <= s_out1(0,2);
	s_in2(59,2) <= s_out2(0,3);

		last_row_cell_3 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,3),
			fetch              => s_fetch(59,3),
			data_in            => s_data_in(59,3),
			data_out           => s_data_out(59,3),
			out1               => s_out1(59,3),
			out2               => s_out2(59,3),
			lock_lower_row_out => s_locks_lower_out(59,3),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,3),
			in2                => s_in2(59,3),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(3)
		);
	s_in1(59,3) <= s_out1(0,3);
	s_in2(59,3) <= s_out2(0,4);

		last_row_cell_4 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,4),
			fetch              => s_fetch(59,4),
			data_in            => s_data_in(59,4),
			data_out           => s_data_out(59,4),
			out1               => s_out1(59,4),
			out2               => s_out2(59,4),
			lock_lower_row_out => s_locks_lower_out(59,4),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,4),
			in2                => s_in2(59,4),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(4)
		);
	s_in1(59,4) <= s_out1(0,4);
	s_in2(59,4) <= s_out2(0,5);

		last_row_cell_5 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,5),
			fetch              => s_fetch(59,5),
			data_in            => s_data_in(59,5),
			data_out           => s_data_out(59,5),
			out1               => s_out1(59,5),
			out2               => s_out2(59,5),
			lock_lower_row_out => s_locks_lower_out(59,5),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,5),
			in2                => s_in2(59,5),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(5)
		);
	s_in1(59,5) <= s_out1(0,5);
	s_in2(59,5) <= s_out2(0,6);

		last_row_cell_6 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,6),
			fetch              => s_fetch(59,6),
			data_in            => s_data_in(59,6),
			data_out           => s_data_out(59,6),
			out1               => s_out1(59,6),
			out2               => s_out2(59,6),
			lock_lower_row_out => s_locks_lower_out(59,6),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,6),
			in2                => s_in2(59,6),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(6)
		);
	s_in1(59,6) <= s_out1(0,6);
	s_in2(59,6) <= s_out2(0,7);

		last_row_cell_7 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,7),
			fetch              => s_fetch(59,7),
			data_in            => s_data_in(59,7),
			data_out           => s_data_out(59,7),
			out1               => s_out1(59,7),
			out2               => s_out2(59,7),
			lock_lower_row_out => s_locks_lower_out(59,7),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,7),
			in2                => s_in2(59,7),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(7)
		);
	s_in1(59,7) <= s_out1(0,7);
	s_in2(59,7) <= s_out2(0,8);

		last_row_cell_8 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,8),
			fetch              => s_fetch(59,8),
			data_in            => s_data_in(59,8),
			data_out           => s_data_out(59,8),
			out1               => s_out1(59,8),
			out2               => s_out2(59,8),
			lock_lower_row_out => s_locks_lower_out(59,8),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,8),
			in2                => s_in2(59,8),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(8)
		);
	s_in1(59,8) <= s_out1(0,8);
	s_in2(59,8) <= s_out2(0,9);

		last_row_cell_9 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,9),
			fetch              => s_fetch(59,9),
			data_in            => s_data_in(59,9),
			data_out           => s_data_out(59,9),
			out1               => s_out1(59,9),
			out2               => s_out2(59,9),
			lock_lower_row_out => s_locks_lower_out(59,9),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,9),
			in2                => s_in2(59,9),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(9)
		);
	s_in1(59,9) <= s_out1(0,9);
	s_in2(59,9) <= s_out2(0,10);

		last_row_cell_10 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,10),
			fetch              => s_fetch(59,10),
			data_in            => s_data_in(59,10),
			data_out           => s_data_out(59,10),
			out1               => s_out1(59,10),
			out2               => s_out2(59,10),
			lock_lower_row_out => s_locks_lower_out(59,10),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,10),
			in2                => s_in2(59,10),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(10)
		);
	s_in1(59,10) <= s_out1(0,10);
	s_in2(59,10) <= s_out2(0,11);

		last_row_cell_11 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,11),
			fetch              => s_fetch(59,11),
			data_in            => s_data_in(59,11),
			data_out           => s_data_out(59,11),
			out1               => s_out1(59,11),
			out2               => s_out2(59,11),
			lock_lower_row_out => s_locks_lower_out(59,11),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,11),
			in2                => s_in2(59,11),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(11)
		);
	s_in1(59,11) <= s_out1(0,11);
	s_in2(59,11) <= s_out2(0,12);

		last_row_cell_12 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,12),
			fetch              => s_fetch(59,12),
			data_in            => s_data_in(59,12),
			data_out           => s_data_out(59,12),
			out1               => s_out1(59,12),
			out2               => s_out2(59,12),
			lock_lower_row_out => s_locks_lower_out(59,12),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,12),
			in2                => s_in2(59,12),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(12)
		);
	s_in1(59,12) <= s_out1(0,12);
	s_in2(59,12) <= s_out2(0,13);

		last_row_cell_13 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,13),
			fetch              => s_fetch(59,13),
			data_in            => s_data_in(59,13),
			data_out           => s_data_out(59,13),
			out1               => s_out1(59,13),
			out2               => s_out2(59,13),
			lock_lower_row_out => s_locks_lower_out(59,13),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,13),
			in2                => s_in2(59,13),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(13)
		);
	s_in1(59,13) <= s_out1(0,13);
	s_in2(59,13) <= s_out2(0,14);

		last_row_cell_14 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,14),
			fetch              => s_fetch(59,14),
			data_in            => s_data_in(59,14),
			data_out           => s_data_out(59,14),
			out1               => s_out1(59,14),
			out2               => s_out2(59,14),
			lock_lower_row_out => s_locks_lower_out(59,14),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,14),
			in2                => s_in2(59,14),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(14)
		);
	s_in1(59,14) <= s_out1(0,14);
	s_in2(59,14) <= s_out2(0,15);

		last_row_cell_15 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,15),
			fetch              => s_fetch(59,15),
			data_in            => s_data_in(59,15),
			data_out           => s_data_out(59,15),
			out1               => s_out1(59,15),
			out2               => s_out2(59,15),
			lock_lower_row_out => s_locks_lower_out(59,15),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,15),
			in2                => s_in2(59,15),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(15)
		);
	s_in1(59,15) <= s_out1(0,15);
	s_in2(59,15) <= s_out2(0,16);

		last_row_cell_16 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,16),
			fetch              => s_fetch(59,16),
			data_in            => s_data_in(59,16),
			data_out           => s_data_out(59,16),
			out1               => s_out1(59,16),
			out2               => s_out2(59,16),
			lock_lower_row_out => s_locks_lower_out(59,16),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,16),
			in2                => s_in2(59,16),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(16)
		);
	s_in1(59,16) <= s_out1(0,16);
	s_in2(59,16) <= s_out2(0,17);

		last_row_cell_17 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,17),
			fetch              => s_fetch(59,17),
			data_in            => s_data_in(59,17),
			data_out           => s_data_out(59,17),
			out1               => s_out1(59,17),
			out2               => s_out2(59,17),
			lock_lower_row_out => s_locks_lower_out(59,17),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,17),
			in2                => s_in2(59,17),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(17)
		);
	s_in1(59,17) <= s_out1(0,17);
	s_in2(59,17) <= s_out2(0,18);

		last_row_cell_18 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,18),
			fetch              => s_fetch(59,18),
			data_in            => s_data_in(59,18),
			data_out           => s_data_out(59,18),
			out1               => s_out1(59,18),
			out2               => s_out2(59,18),
			lock_lower_row_out => s_locks_lower_out(59,18),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,18),
			in2                => s_in2(59,18),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(18)
		);
	s_in1(59,18) <= s_out1(0,18);
	s_in2(59,18) <= s_out2(0,19);

		last_row_cell_19 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,19),
			fetch              => s_fetch(59,19),
			data_in            => s_data_in(59,19),
			data_out           => s_data_out(59,19),
			out1               => s_out1(59,19),
			out2               => s_out2(59,19),
			lock_lower_row_out => s_locks_lower_out(59,19),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,19),
			in2                => s_in2(59,19),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(19)
		);
	s_in1(59,19) <= s_out1(0,19);
	s_in2(59,19) <= s_out2(0,20);

		last_row_cell_20 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,20),
			fetch              => s_fetch(59,20),
			data_in            => s_data_in(59,20),
			data_out           => s_data_out(59,20),
			out1               => s_out1(59,20),
			out2               => s_out2(59,20),
			lock_lower_row_out => s_locks_lower_out(59,20),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,20),
			in2                => s_in2(59,20),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(20)
		);
	s_in1(59,20) <= s_out1(0,20);
	s_in2(59,20) <= s_out2(0,21);

		last_row_cell_21 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,21),
			fetch              => s_fetch(59,21),
			data_in            => s_data_in(59,21),
			data_out           => s_data_out(59,21),
			out1               => s_out1(59,21),
			out2               => s_out2(59,21),
			lock_lower_row_out => s_locks_lower_out(59,21),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,21),
			in2                => s_in2(59,21),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(21)
		);
	s_in1(59,21) <= s_out1(0,21);
	s_in2(59,21) <= s_out2(0,22);

		last_row_cell_22 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,22),
			fetch              => s_fetch(59,22),
			data_in            => s_data_in(59,22),
			data_out           => s_data_out(59,22),
			out1               => s_out1(59,22),
			out2               => s_out2(59,22),
			lock_lower_row_out => s_locks_lower_out(59,22),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,22),
			in2                => s_in2(59,22),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(22)
		);
	s_in1(59,22) <= s_out1(0,22);
	s_in2(59,22) <= s_out2(0,23);

		last_row_cell_23 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,23),
			fetch              => s_fetch(59,23),
			data_in            => s_data_in(59,23),
			data_out           => s_data_out(59,23),
			out1               => s_out1(59,23),
			out2               => s_out2(59,23),
			lock_lower_row_out => s_locks_lower_out(59,23),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,23),
			in2                => s_in2(59,23),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(23)
		);
	s_in1(59,23) <= s_out1(0,23);
	s_in2(59,23) <= s_out2(0,24);

		last_row_cell_24 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,24),
			fetch              => s_fetch(59,24),
			data_in            => s_data_in(59,24),
			data_out           => s_data_out(59,24),
			out1               => s_out1(59,24),
			out2               => s_out2(59,24),
			lock_lower_row_out => s_locks_lower_out(59,24),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,24),
			in2                => s_in2(59,24),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(24)
		);
	s_in1(59,24) <= s_out1(0,24);
	s_in2(59,24) <= s_out2(0,25);

		last_row_cell_25 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,25),
			fetch              => s_fetch(59,25),
			data_in            => s_data_in(59,25),
			data_out           => s_data_out(59,25),
			out1               => s_out1(59,25),
			out2               => s_out2(59,25),
			lock_lower_row_out => s_locks_lower_out(59,25),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,25),
			in2                => s_in2(59,25),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(25)
		);
	s_in1(59,25) <= s_out1(0,25);
	s_in2(59,25) <= s_out2(0,26);

		last_row_cell_26 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,26),
			fetch              => s_fetch(59,26),
			data_in            => s_data_in(59,26),
			data_out           => s_data_out(59,26),
			out1               => s_out1(59,26),
			out2               => s_out2(59,26),
			lock_lower_row_out => s_locks_lower_out(59,26),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,26),
			in2                => s_in2(59,26),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(26)
		);
	s_in1(59,26) <= s_out1(0,26);
	s_in2(59,26) <= s_out2(0,27);

		last_row_cell_27 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,27),
			fetch              => s_fetch(59,27),
			data_in            => s_data_in(59,27),
			data_out           => s_data_out(59,27),
			out1               => s_out1(59,27),
			out2               => s_out2(59,27),
			lock_lower_row_out => s_locks_lower_out(59,27),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,27),
			in2                => s_in2(59,27),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(27)
		);
	s_in1(59,27) <= s_out1(0,27);
	s_in2(59,27) <= s_out2(0,28);

		last_row_cell_28 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,28),
			fetch              => s_fetch(59,28),
			data_in            => s_data_in(59,28),
			data_out           => s_data_out(59,28),
			out1               => s_out1(59,28),
			out2               => s_out2(59,28),
			lock_lower_row_out => s_locks_lower_out(59,28),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,28),
			in2                => s_in2(59,28),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(28)
		);
	s_in1(59,28) <= s_out1(0,28);
	s_in2(59,28) <= s_out2(0,29);

		last_row_cell_29 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,29),
			fetch              => s_fetch(59,29),
			data_in            => s_data_in(59,29),
			data_out           => s_data_out(59,29),
			out1               => s_out1(59,29),
			out2               => s_out2(59,29),
			lock_lower_row_out => s_locks_lower_out(59,29),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,29),
			in2                => s_in2(59,29),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(29)
		);
	s_in1(59,29) <= s_out1(0,29);
	s_in2(59,29) <= s_out2(0,30);

		last_row_cell_30 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,30),
			fetch              => s_fetch(59,30),
			data_in            => s_data_in(59,30),
			data_out           => s_data_out(59,30),
			out1               => s_out1(59,30),
			out2               => s_out2(59,30),
			lock_lower_row_out => s_locks_lower_out(59,30),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,30),
			in2                => s_in2(59,30),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(30)
		);
	s_in1(59,30) <= s_out1(0,30);
	s_in2(59,30) <= s_out2(0,31);

		last_row_cell_31 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,31),
			fetch              => s_fetch(59,31),
			data_in            => s_data_in(59,31),
			data_out           => s_data_out(59,31),
			out1               => s_out1(59,31),
			out2               => s_out2(59,31),
			lock_lower_row_out => s_locks_lower_out(59,31),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,31),
			in2                => s_in2(59,31),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(31)
		);
	s_in1(59,31) <= s_out1(0,31);
	s_in2(59,31) <= s_out2(0,32);

		last_row_cell_32 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,32),
			fetch              => s_fetch(59,32),
			data_in            => s_data_in(59,32),
			data_out           => s_data_out(59,32),
			out1               => s_out1(59,32),
			out2               => s_out2(59,32),
			lock_lower_row_out => s_locks_lower_out(59,32),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,32),
			in2                => s_in2(59,32),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(32)
		);
	s_in1(59,32) <= s_out1(0,32);
	s_in2(59,32) <= s_out2(0,33);

		last_row_cell_33 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,33),
			fetch              => s_fetch(59,33),
			data_in            => s_data_in(59,33),
			data_out           => s_data_out(59,33),
			out1               => s_out1(59,33),
			out2               => s_out2(59,33),
			lock_lower_row_out => s_locks_lower_out(59,33),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,33),
			in2                => s_in2(59,33),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(33)
		);
	s_in1(59,33) <= s_out1(0,33);
	s_in2(59,33) <= s_out2(0,34);

		last_row_cell_34 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,34),
			fetch              => s_fetch(59,34),
			data_in            => s_data_in(59,34),
			data_out           => s_data_out(59,34),
			out1               => s_out1(59,34),
			out2               => s_out2(59,34),
			lock_lower_row_out => s_locks_lower_out(59,34),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,34),
			in2                => s_in2(59,34),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(34)
		);
	s_in1(59,34) <= s_out1(0,34);
	s_in2(59,34) <= s_out2(0,35);

		last_row_cell_35 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,35),
			fetch              => s_fetch(59,35),
			data_in            => s_data_in(59,35),
			data_out           => s_data_out(59,35),
			out1               => s_out1(59,35),
			out2               => s_out2(59,35),
			lock_lower_row_out => s_locks_lower_out(59,35),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,35),
			in2                => s_in2(59,35),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(35)
		);
	s_in1(59,35) <= s_out1(0,35);
	s_in2(59,35) <= s_out2(0,36);

		last_row_cell_36 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,36),
			fetch              => s_fetch(59,36),
			data_in            => s_data_in(59,36),
			data_out           => s_data_out(59,36),
			out1               => s_out1(59,36),
			out2               => s_out2(59,36),
			lock_lower_row_out => s_locks_lower_out(59,36),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,36),
			in2                => s_in2(59,36),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(36)
		);
	s_in1(59,36) <= s_out1(0,36);
	s_in2(59,36) <= s_out2(0,37);

		last_row_cell_37 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,37),
			fetch              => s_fetch(59,37),
			data_in            => s_data_in(59,37),
			data_out           => s_data_out(59,37),
			out1               => s_out1(59,37),
			out2               => s_out2(59,37),
			lock_lower_row_out => s_locks_lower_out(59,37),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,37),
			in2                => s_in2(59,37),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(37)
		);
	s_in1(59,37) <= s_out1(0,37);
	s_in2(59,37) <= s_out2(0,38);

		last_row_cell_38 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,38),
			fetch              => s_fetch(59,38),
			data_in            => s_data_in(59,38),
			data_out           => s_data_out(59,38),
			out1               => s_out1(59,38),
			out2               => s_out2(59,38),
			lock_lower_row_out => s_locks_lower_out(59,38),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,38),
			in2                => s_in2(59,38),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(38)
		);
	s_in1(59,38) <= s_out1(0,38);
	s_in2(59,38) <= s_out2(0,39);

		last_row_cell_39 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,39),
			fetch              => s_fetch(59,39),
			data_in            => s_data_in(59,39),
			data_out           => s_data_out(59,39),
			out1               => s_out1(59,39),
			out2               => s_out2(59,39),
			lock_lower_row_out => s_locks_lower_out(59,39),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,39),
			in2                => s_in2(59,39),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(39)
		);
	s_in1(59,39) <= s_out1(0,39);
	s_in2(59,39) <= s_out2(0,40);

		last_row_cell_40 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,40),
			fetch              => s_fetch(59,40),
			data_in            => s_data_in(59,40),
			data_out           => s_data_out(59,40),
			out1               => s_out1(59,40),
			out2               => s_out2(59,40),
			lock_lower_row_out => s_locks_lower_out(59,40),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,40),
			in2                => s_in2(59,40),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(40)
		);
	s_in1(59,40) <= s_out1(0,40);
	s_in2(59,40) <= s_out2(0,41);

		last_row_cell_41 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,41),
			fetch              => s_fetch(59,41),
			data_in            => s_data_in(59,41),
			data_out           => s_data_out(59,41),
			out1               => s_out1(59,41),
			out2               => s_out2(59,41),
			lock_lower_row_out => s_locks_lower_out(59,41),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,41),
			in2                => s_in2(59,41),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(41)
		);
	s_in1(59,41) <= s_out1(0,41);
	s_in2(59,41) <= s_out2(0,42);

		last_row_cell_42 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,42),
			fetch              => s_fetch(59,42),
			data_in            => s_data_in(59,42),
			data_out           => s_data_out(59,42),
			out1               => s_out1(59,42),
			out2               => s_out2(59,42),
			lock_lower_row_out => s_locks_lower_out(59,42),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,42),
			in2                => s_in2(59,42),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(42)
		);
	s_in1(59,42) <= s_out1(0,42);
	s_in2(59,42) <= s_out2(0,43);

		last_row_cell_43 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,43),
			fetch              => s_fetch(59,43),
			data_in            => s_data_in(59,43),
			data_out           => s_data_out(59,43),
			out1               => s_out1(59,43),
			out2               => s_out2(59,43),
			lock_lower_row_out => s_locks_lower_out(59,43),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,43),
			in2                => s_in2(59,43),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(43)
		);
	s_in1(59,43) <= s_out1(0,43);
	s_in2(59,43) <= s_out2(0,44);

		last_row_cell_44 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,44),
			fetch              => s_fetch(59,44),
			data_in            => s_data_in(59,44),
			data_out           => s_data_out(59,44),
			out1               => s_out1(59,44),
			out2               => s_out2(59,44),
			lock_lower_row_out => s_locks_lower_out(59,44),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,44),
			in2                => s_in2(59,44),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(44)
		);
	s_in1(59,44) <= s_out1(0,44);
	s_in2(59,44) <= s_out2(0,45);

		last_row_cell_45 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,45),
			fetch              => s_fetch(59,45),
			data_in            => s_data_in(59,45),
			data_out           => s_data_out(59,45),
			out1               => s_out1(59,45),
			out2               => s_out2(59,45),
			lock_lower_row_out => s_locks_lower_out(59,45),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,45),
			in2                => s_in2(59,45),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(45)
		);
	s_in1(59,45) <= s_out1(0,45);
	s_in2(59,45) <= s_out2(0,46);

		last_row_cell_46 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,46),
			fetch              => s_fetch(59,46),
			data_in            => s_data_in(59,46),
			data_out           => s_data_out(59,46),
			out1               => s_out1(59,46),
			out2               => s_out2(59,46),
			lock_lower_row_out => s_locks_lower_out(59,46),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,46),
			in2                => s_in2(59,46),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(46)
		);
	s_in1(59,46) <= s_out1(0,46);
	s_in2(59,46) <= s_out2(0,47);

		last_row_cell_47 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,47),
			fetch              => s_fetch(59,47),
			data_in            => s_data_in(59,47),
			data_out           => s_data_out(59,47),
			out1               => s_out1(59,47),
			out2               => s_out2(59,47),
			lock_lower_row_out => s_locks_lower_out(59,47),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,47),
			in2                => s_in2(59,47),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(47)
		);
	s_in1(59,47) <= s_out1(0,47);
	s_in2(59,47) <= s_out2(0,48);

		last_row_cell_48 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,48),
			fetch              => s_fetch(59,48),
			data_in            => s_data_in(59,48),
			data_out           => s_data_out(59,48),
			out1               => s_out1(59,48),
			out2               => s_out2(59,48),
			lock_lower_row_out => s_locks_lower_out(59,48),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,48),
			in2                => s_in2(59,48),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(48)
		);
	s_in1(59,48) <= s_out1(0,48);
	s_in2(59,48) <= s_out2(0,49);

		last_row_cell_49 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,49),
			fetch              => s_fetch(59,49),
			data_in            => s_data_in(59,49),
			data_out           => s_data_out(59,49),
			out1               => s_out1(59,49),
			out2               => s_out2(59,49),
			lock_lower_row_out => s_locks_lower_out(59,49),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,49),
			in2                => s_in2(59,49),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(49)
		);
	s_in1(59,49) <= s_out1(0,49);
	s_in2(59,49) <= s_out2(0,50);

		last_row_cell_50 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,50),
			fetch              => s_fetch(59,50),
			data_in            => s_data_in(59,50),
			data_out           => s_data_out(59,50),
			out1               => s_out1(59,50),
			out2               => s_out2(59,50),
			lock_lower_row_out => s_locks_lower_out(59,50),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,50),
			in2                => s_in2(59,50),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(50)
		);
	s_in1(59,50) <= s_out1(0,50);
	s_in2(59,50) <= s_out2(0,51);

		last_row_cell_51 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,51),
			fetch              => s_fetch(59,51),
			data_in            => s_data_in(59,51),
			data_out           => s_data_out(59,51),
			out1               => s_out1(59,51),
			out2               => s_out2(59,51),
			lock_lower_row_out => s_locks_lower_out(59,51),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,51),
			in2                => s_in2(59,51),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(51)
		);
	s_in1(59,51) <= s_out1(0,51);
	s_in2(59,51) <= s_out2(0,52);

		last_row_cell_52 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,52),
			fetch              => s_fetch(59,52),
			data_in            => s_data_in(59,52),
			data_out           => s_data_out(59,52),
			out1               => s_out1(59,52),
			out2               => s_out2(59,52),
			lock_lower_row_out => s_locks_lower_out(59,52),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,52),
			in2                => s_in2(59,52),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(52)
		);
	s_in1(59,52) <= s_out1(0,52);
	s_in2(59,52) <= s_out2(0,53);

		last_row_cell_53 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,53),
			fetch              => s_fetch(59,53),
			data_in            => s_data_in(59,53),
			data_out           => s_data_out(59,53),
			out1               => s_out1(59,53),
			out2               => s_out2(59,53),
			lock_lower_row_out => s_locks_lower_out(59,53),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,53),
			in2                => s_in2(59,53),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(53)
		);
	s_in1(59,53) <= s_out1(0,53);
	s_in2(59,53) <= s_out2(0,54);

		last_row_cell_54 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,54),
			fetch              => s_fetch(59,54),
			data_in            => s_data_in(59,54),
			data_out           => s_data_out(59,54),
			out1               => s_out1(59,54),
			out2               => s_out2(59,54),
			lock_lower_row_out => s_locks_lower_out(59,54),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,54),
			in2                => s_in2(59,54),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(54)
		);
	s_in1(59,54) <= s_out1(0,54);
	s_in2(59,54) <= s_out2(0,55);

		last_row_cell_55 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,55),
			fetch              => s_fetch(59,55),
			data_in            => s_data_in(59,55),
			data_out           => s_data_out(59,55),
			out1               => s_out1(59,55),
			out2               => s_out2(59,55),
			lock_lower_row_out => s_locks_lower_out(59,55),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,55),
			in2                => s_in2(59,55),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(55)
		);
	s_in1(59,55) <= s_out1(0,55);
	s_in2(59,55) <= s_out2(0,56);

		last_row_cell_56 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,56),
			fetch              => s_fetch(59,56),
			data_in            => s_data_in(59,56),
			data_out           => s_data_out(59,56),
			out1               => s_out1(59,56),
			out2               => s_out2(59,56),
			lock_lower_row_out => s_locks_lower_out(59,56),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,56),
			in2                => s_in2(59,56),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(56)
		);
	s_in1(59,56) <= s_out1(0,56);
	s_in2(59,56) <= s_out2(0,57);

		last_row_cell_57 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,57),
			fetch              => s_fetch(59,57),
			data_in            => s_data_in(59,57),
			data_out           => s_data_out(59,57),
			out1               => s_out1(59,57),
			out2               => s_out2(59,57),
			lock_lower_row_out => s_locks_lower_out(59,57),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,57),
			in2                => s_in2(59,57),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(57)
		);
	s_in1(59,57) <= s_out1(0,57);
	s_in2(59,57) <= s_out2(0,58);

		last_row_cell_58 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,58),
			fetch              => s_fetch(59,58),
			data_in            => s_data_in(59,58),
			data_out           => s_data_out(59,58),
			out1               => s_out1(59,58),
			out2               => s_out2(59,58),
			lock_lower_row_out => s_locks_lower_out(59,58),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,58),
			in2                => s_in2(59,58),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(58)
		);
	s_in1(59,58) <= s_out1(0,58);
	s_in2(59,58) <= s_out2(0,59);

		last_row_cell_59 : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,59),
			fetch              => s_fetch(59,59),
			data_in            => s_data_in(59,59),
			data_out           => s_data_out(59,59),
			out1               => s_out1(59,59),
			out2               => s_out2(59,59),
			lock_lower_row_out => s_locks_lower_out(59,59),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,59),
			in2                => s_in2(59,59),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(59)
		);
	s_in1(59,59) <= s_out1(0,59);
	s_in2(59,59) <= s_out2(0,60);

		last_cell : basic_cell port map(
			clk                => clk,
			rst                => rst,
			en                 => en,
			load               => s_load(59,60),
			fetch              => s_fetch(59,60),
			data_in            => s_data_in(59,60),
			data_out           => s_data_out(59,60),
			out1               => s_out1(59,60),
			out2               => s_out2(59,60),
			lock_lower_row_out => s_locks_lower_out(59,60),
			lock_lower_row_in  => '0',
			in1                => s_in1(59,60),
			in2                => (others => '0'),
			lock_row           => s_locks(59),
			piv_found          => s_piv_found,
			row_data           => s_row_data(59),
			col_data           => s_col_data(60)
		);
	s_in1(59,60) <= s_out1(0,60);

	en   <= enable;
	done <= check_locks(s_locks);

	process(clk)
		variable v_i : integer range 0 to ROWS-1;
		variable v_j : integer range 0 to COLS-1;
	begin
		if (rising_edge(clk)) then
			if (rst = '1') then
				v_i := 0;
				v_j := 0;
				
			else
				v_i := to_integer(unsigned(i));
				v_j := to_integer(unsigned(j));

				if (lo = '1') then
					s_load(v_i,v_j)    <= '1';
					s_data_in(v_i,v_j) <= data_in;
				else
					s_load(v_i,v_j) <= '0';
				end if;

				if(fet = '1') then
					s_fetch(v_i,v_j) <= '1';
					data_out         <= s_data_out(v_i,v_j);
				else
					s_fetch(v_i,v_j) <= '0';
				end if;
			end if;
		end if;
	end process;
end architecture behav;
